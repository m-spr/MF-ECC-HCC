LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity top_module_for_mem_free_ECC_10000 is
    generic (
        dimension_size     : integer := 10240;   -- dimension size 
        dimension_WIDTH    : integer := 14;     -- log2 dimension size 
        dimension_segmentation    : integer := 1280;     -- genrate input
        class_size    : integer := 10;     -- number of classes
        ECC_WIDTH          : integer := 5       -- bit-width of ECC_code 
    );
    port (
	clk                     : in std_logic;
    rst                     : in std_logic;
    pop_en                  : in std_logic;
	din 					: in std_logic_vector((dimension_size/dimension_segmentation)-1 downto 0);
    count_sim     :out std_logic_vector(dimension_WIDTH-1 downto 0)
	);	
end entity;

architecture behavior of top_module_for_mem_free_ECC_10000 is

component reading_normal is
    generic (
        dimension_size     : integer := 1024;   -- dimension size 
        dimension_WIDTH    : integer := 10;     -- log2 dimension size 
        class_size    : integer := 10;     -- number of classes
        ECC_WIDTH          : integer := 8       -- bit-width of ECC_code 
    );
	port (
	clk                     : in std_logic;
    rst                     : in std_logic;
	din 					: in std_logic_vector(dimension_size-1 downto 0);
    count_reg               : in std_logic_vector(dimension_WIDTH-1 downto 0);
    dout                    : out std_logic_vector(dimension_WIDTH-1 downto 0)
	);	
end component;



component popCount IS
	GENERIC (lenPop : INTEGER := 8);   -- bit width out popCounters --- LOG2(#feature)
	PORT (
		clk , rst 	: IN STD_LOGIC;
		en		 	: IN STD_LOGIC;
		dout        : OUT  STD_LOGIC_VECTOR (lenPop-1 DOWNTO 0)
	);
END component;


signal realdin 					:  std_logic_vector((dimension_size)-1 downto 0);

type index_array is array (0 to dimension_size-1) of std_logic_vector(dimension_WIDTH-1 downto 0);
    
signal index_memory               : index_array;
signal count_reg               :  std_logic_vector(dimension_WIDTH-1 downto 0);
       
begin

    input_gen: for k in 0 to dimension_segmentation-1 generate
        realdin((dimension_size/dimension_segmentation)*(k+1)-1 downto (dimension_size/dimension_segmentation)*k) <= din;
    end generate;
    
    
    ECCuutMem: entity work.reading_normal 
	generic map(
		dimension_size  => dimension_size,
        dimension_WIDTH  => dimension_WIDTH,
        class_size  =>  class_size,
        ECC_WIDTH => ECC_WIDTH)
	port map(
		clk  => clk,
		rst  => rst,
		din  => realdin,
	    count_reg 		=> count_reg,
		dout  => count_sim
		);

    -- Count_reg counter
    counter: entity work.popCount 
        generic map(lenPop => dimension_WIDTH)
        port map(
            clk  => clk,
            rst  => rst,
            en   => pop_en,
            dout => count_reg
        );

end architecture;


----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ECC_vhdl_module is
    generic (
        C      : integer := 10;        -- Bit width number of classes or the segments size that we are going to correct
        ECC_bit: integer := 5          -- Number of bits for correction each column
    );
    port (
        d           : in  std_logic_vector(C-1 downto 0);  -- Input data vector
        p           : in  std_logic_vector(ECC_bit-1 downto 0);  -- Input ECC bits
        double_error: out std_logic;                        -- Output flag for double error
        dcw         : out std_logic_vector(C-1 downto 0)    -- Corrected data vector
    );
end entity ECC_vhdl_module;

architecture Behavioral of ECC_vhdl_module is
    signal dp : std_logic_vector(4 downto 0);  -- Parity calculated from input data
    signal s  : std_logic_vector(4 downto 0);  -- Syndrome bits
    signal df : std_logic_vector(9 downto 0);  -- Flag bit for getting correct data
    signal xw : std_logic;                     -- Intermediate signal for double error flag
begin

    -- Data Parity calculation
    dp(0) <= d(0) xor d(1) xor d(3) xor d(4) xor d(6) xor d(8);
    dp(1) <= d(0) xor d(2) xor d(3) xor d(5) xor d(6) xor d(9);
    dp(2) <= d(1) xor d(2) xor d(3) xor d(7) xor d(8) xor d(9);
    dp(3) <= d(4) xor d(5) xor d(6) xor d(7) xor d(8) xor d(9);
    dp(4) <= d(0) xor d(1) xor d(2) xor d(3) xor d(4) xor d(5) xor d(6) xor d(7) xor d(8) xor d(9) xor p(0) xor p(1) xor p(2) xor p(3);

    -- Syndrome: xor with actual parity
    s(0) <= p(0) xor dp(0);
    s(1) <= p(1) xor dp(1);
    s(2) <= p(2) xor dp(2);
    s(3) <= p(3) xor dp(3);
    s(4) <= p(4) xor dp(4);

    -- Flag bit for getting correct data
    df(0) <= s(0) and s(1) and not s(2) and not s(3) and s(4);
    df(1) <= s(0) and not s(1) and s(2) and not s(3) and s(4);
    df(2) <= not s(0) and s(1) and s(2) and not s(3) and s(4);
    df(3) <= s(0) and s(1) and s(2) and not s(3) and s(4);
    df(4) <= s(0) and not s(1) and not s(2) and s(3) and s(4);
    df(5) <= not s(0) and s(1) and not s(2) and s(3) and s(4);
    df(6) <= s(0) and s(1) and not s(2) and s(3) and s(4);
    df(7) <= not s(0) and not s(1) and s(2) and s(3) and s(4);
    df(8) <= s(0) and not s(1) and s(2) and s(3) and s(4);
    df(9) <= not s(0) and s(1) and s(2) and s(3) and s(4);

    -- Corrected data bits
    dcw(0) <= df(0) xor d(0);
    dcw(1) <= df(1) xor d(1);
    dcw(2) <= df(2) xor d(2);
    dcw(3) <= df(3) xor d(3);
    dcw(4) <= df(4) xor d(4);
    dcw(5) <= df(5) xor d(5);
    dcw(6) <= df(6) xor d(6);
    dcw(7) <= df(7) xor d(7);
    dcw(8) <= df(8) xor d(8);
    dcw(9) <= df(9) xor d(9);

    -- Intermediate signal for double error flag
    xw <= s(0) or s(1) or s(2) or s(3);

    -- Flag for double error
    double_error <= not s(4) and xw;  -- If 1, that means double error exists

end architecture Behavioral;


---------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY popCount IS
	GENERIC (lenPop : INTEGER := 8);   -- bit width out popCounters --- LOG2(#feature)
	PORT (
		clk , rst 	: IN STD_LOGIC;
		en		 	: IN STD_LOGIC;
		dout        : OUT  STD_LOGIC_VECTOR (lenPop-1 DOWNTO 0)
	);
END ENTITY popCount;

ARCHITECTURE behavioral OF popCount IS
SIGNAL popOut : STD_LOGIC_VECTOR (lenPop - 1 DOWNTO 0);
	
BEGIN

	PROCESS(clk)
		BEGIN 
		    IF rising_edge(clk) THEN
			    IF(rst = '1')THEN
				   popOut <= (OTHERS=>'0');
				ELSIF (en ='1') THEN 
				   popOut <= STD_LOGIC_VECTOR (UNSIGNED(popOut) + 1);
				END IF;
			END IF;
	END PROCESS;

	dout <= popOut;
END ARCHITECTURE behavioral;

---------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CHV_mem_10000 is
    Port (
        clk     : in  STD_LOGIC;
        address : in  STD_LOGIC_VECTOR(13 downto 0);
        data    : out STD_LOGIC_VECTOR(10 downto 0)
    );
end CHV_mem_10000;

architecture Behavioral of CHV_mem_10000 is
begin
    process(clk)
    begin
        if rising_edge(clk) then
            case address is
                when x"00" => data <= "1010110001";
                when x"01" => data <= "0100000000";
                when x"02" => data <= "0010101000";
                when x"03" => data <= "0100000000";
                when x"04" => data <= "1001010000";
                when x"05" => data <= "1011011011";
                when x"06" => data <= "0100000000";
                when x"07" => data <= "0100000000";
                when x"08" => data <= "0100000000";
                when x"09" => data <= "0010101000";
                when x"0A" => data <= "1110100111";
                when x"0B" => data <= "0100000000";
                when x"0C" => data <= "0100000000";
                when x"0D" => data <= "1001010000";
                when x"0E" => data <= "0100000000";
                when x"0F" => data <= "0100000000";
                when x"10" => data <= "0100110101";
                when x"11" => data <= "1111111000";
                when x"12" => data <= "1001010000";
                when x"13" => data <= "0100000000";
                when x"14" => data <= "1010000100";
                when x"15" => data <= "1011011011";
                when x"16" => data <= "0100000000";
                when x"17" => data <= "0100000000";
                when x"18" => data <= "0100000000";
                when x"19" => data <= "0100000000";
                when x"1A" => data <= "0100000000";
                when x"1B" => data <= "0011000010";
                when x"1C" => data <= "0100000000";
                when x"1D" => data <= "1001010000";
                when x"1E" => data <= "0100000000";
                when x"1F" => data <= "1000111010";
                when x"20" => data <= "0100000000";
                when x"21" => data <= "0100000000";
                when x"22" => data <= "0000100011";
                when x"23" => data <= "0100000000";
                when x"24" => data <= "0100000000";
                when x"25" => data <= "0100000000";
                when x"26" => data <= "1001010000";
                when x"27" => data <= "0100000000";
                when x"28" => data <= "0100000000";
                when x"29" => data <= "0100000000";
                when x"2A" => data <= "0100000000";
                when x"2B" => data <= "0100000000";
                when x"2C" => data <= "1001010000";
                when x"2D" => data <= "0100110101";
                when x"2E" => data <= "0100000000";
                when x"2F" => data <= "0100000000";
                when x"30" => data <= "0100000000";
                when x"31" => data <= "0100000000";
                when x"32" => data <= "0011000010";
                when x"33" => data <= "0100000000";
                when x"34" => data <= "0100000000";
                when x"35" => data <= "1001010000";
                when x"36" => data <= "0100000000";
                when x"37" => data <= "1001010000";
                when x"38" => data <= "0101011111";
                when x"39" => data <= "1001010000";
                when x"3A" => data <= "0100000000";
                when x"3B" => data <= "0110001011";
                when x"3C" => data <= "0100000000";
                when x"3D" => data <= "1110010010";
                when x"3E" => data <= "0100000000";
                when x"3F" => data <= "0101011111";
                when x"40" => data <= "0100000000";
                when x"41" => data <= "1010000100";
                when x"42" => data <= "0100000000";
                when x"43" => data <= "1111001101";
                when x"44" => data <= "0100000000";
                when x"45" => data <= "0100000000";
                when x"46" => data <= "0100000000";
                when x"47" => data <= "0100000000";
                when x"48" => data <= "0100110101";
                when x"49" => data <= "0100000000";
                when x"4A" => data <= "0011000010";
                when x"4B" => data <= "0100000000";
                when x"4C" => data <= "0100000000";
                when x"4D" => data <= "0100000000";
                when x"4E" => data <= "1101000110";
                when x"4F" => data <= "0100000000";
                when x"50" => data <= "1001010000";
                when x"51" => data <= "0100110101";
                when x"52" => data <= "0100000000";
                when x"53" => data <= "0100000000";
                when x"54" => data <= "0111100001";
                when x"55" => data <= "0100000000";
                when x"56" => data <= "1001010000";
                when x"57" => data <= "0100000000";
                when x"58" => data <= "0100000000";
                when x"59" => data <= "1110100111";
                when x"5A" => data <= "0100000000";
                when x"5B" => data <= "0010101000";
                when x"5C" => data <= "0100000000";
                when x"5D" => data <= "0100000000";
                when x"5E" => data <= "0100110101";
                when x"5F" => data <= "0100110101";
                when x"60" => data <= "0100000000";
                when x"61" => data <= "0100000000";
                when x"62" => data <= "0100000000";
                when x"63" => data <= "0100000000";
                when x"64" => data <= "1111111000";
                when x"65" => data <= "0010101000";
                when x"66" => data <= "0100000000";
                when x"67" => data <= "0100000000";
                when x"68" => data <= "0101011111";
                when x"69" => data <= "0010101000";
                when x"6A" => data <= "1111111000";
                when x"6B" => data <= "0100000000";
                when x"6C" => data <= "1001111111";
                when x"6D" => data <= "1000010101";
                when x"6E" => data <= "1111010111";
                when x"6F" => data <= "0111111011";
                when x"70" => data <= "1001111111";
                when x"71" => data <= "0111001110";
                when x"72" => data <= "1010101011";
                when x"73" => data <= "1110111101";
                when x"74" => data <= "0111111011";
                when x"75" => data <= "0101110000";
                when x"76" => data <= "1001111111";
                when x"77" => data <= "1111010111";
                when x"78" => data <= "0111111011";
                when x"79" => data <= "1001111111";
                when x"7A" => data <= "0000001100";
                when x"7B" => data <= "0101110000";
                when x"7C" => data <= "1000100000";
                when x"7D" => data <= "1001111111";
                when x"7E" => data <= "1001111111";
                when x"7F" => data <= "1110111101";
                when x"80" => data <= "1111010111";
                when x"81" => data <= "1110111101";
                when x"82" => data <= "0111111011";
                when x"83" => data <= "0011101101";
                when x"84" => data <= "0101000101";
                when x"85" => data <= "0111111011";
                when x"86" => data <= "0100101111";
                when x"87" => data <= "0100101111";
                when x"88" => data <= "0111111011";
                when x"89" => data <= "1110001000";
                when x"8A" => data <= "0100101111";
                when x"8B" => data <= "1111010111";
                when x"8C" => data <= "1001111111";
                when x"8D" => data <= "1111010111";
                when x"8E" => data <= "0111111011";
                when x"8F" => data <= "1001111111";
                when x"90" => data <= "0111111011";
                when x"91" => data <= "1110111101";
                when x"92" => data <= "1000100000";
                when x"93" => data <= "0001010011";
                when x"94" => data <= "1001111111";
                when x"95" => data <= "0111001110";
                when x"96" => data <= "0111111011";
                when x"97" => data <= "0111111011";
                when x"98" => data <= "1001111111";
                when x"99" => data <= "0111111011";
                when x"9A" => data <= "0111111011";
                when x"9B" => data <= "0111001110";
                when x"9C" => data <= "0000001100";
                when x"9D" => data <= "0101000101";
                when x"9E" => data <= "1110111101";
                when x"9F" => data <= "0111111011";
                when x"A0" => data <= "1000010101";
                when x"A1" => data <= "1110001000";
                when x"A2" => data <= "1101011100";
                when x"A3" => data <= "1001111111";
                when x"A4" => data <= "0011011000";
                when x"A5" => data <= "1110001000";
                when x"A6" => data <= "1110111101";
                when x"A7" => data <= "0101000101";
                when x"A8" => data <= "0100101111";
                when x"A9" => data <= "0111001110";
                when x"AA" => data <= "1110111101";
                when x"AB" => data <= "0110000110";
                when x"AC" => data <= "1100010100";
                when x"AD" => data <= "0101010010";
                when x"AE" => data <= "1111000000";
                when x"AF" => data <= "1000000010";
                when x"B0" => data <= "0110000110";
                when x"B1" => data <= "1111110101";
                when x"B2" => data <= "1111000000";
                when x"B3" => data <= "0001000100";
                when x"B4" => data <= "0100111000";
                when x"B5" => data <= "0001000100";
                when x"B6" => data <= "1000110111";
                when x"B7" => data <= "1111110101";
                when x"B8" => data <= "1011010110";
                when x"B9" => data <= "0100001101";
                when x"BA" => data <= "0001000100";
                when x"BB" => data <= "0001000100";
                when x"BC" => data <= "0100001101";
                when x"BD" => data <= "1111000000";
                when x"BE" => data <= "0100111000";
                when x"BF" => data <= "1000110111";
                when x"C0" => data <= "1011100011";
                when x"C1" => data <= "1111000000";
                when x"C2" => data <= "0101010010";
                when x"C3" => data <= "1111000000";
                when x"C4" => data <= "1111110101";
                when x"C5" => data <= "0001000100";
                when x"C6" => data <= "0101010010";
                when x"C7" => data <= "1001011101";
                when x"C8" => data <= "0001000100";
                when x"C9" => data <= "1000000010";
                when x"CA" => data <= "0001000100";
                when x"CB" => data <= "0011111010";
                when x"CC" => data <= "0100001101";
                when x"CD" => data <= "0001000100";
                when x"CE" => data <= "0101100111";
                when x"CF" => data <= "1100010100";
                when x"D0" => data <= "0101010010";
                when x"D1" => data <= "0110000110";
                when x"D2" => data <= "0010100101";
                when x"D3" => data <= "1111011010";
                when x"D4" => data <= "1111011010";
                when x"D5" => data <= "1111011010";
                when x"D6" => data <= "1001110010";
                when x"D7" => data <= "0101001000";
                when x"D8" => data <= "0000000001";
                when x"D9" => data <= "1111101111";
                when x"DA" => data <= "1111011010";
                when x"DB" => data <= "1111011010";
                when x"DC" => data <= "1111101111";
                when x"DD" => data <= "1111011010";
                when x"DE" => data <= "1011001100";
                when x"DF" => data <= "1000011000";
                when x"E0" => data <= "0010111111";
                when x"E1" => data <= "1111101111";
                when x"E2" => data <= "1011111001";
                when x"E3" => data <= "1111101111";
                when x"E4" => data <= "1111011010";
                when x"E5" => data <= "1111011010";
                when x"E6" => data <= "1111011010";
                when x"E7" => data <= "1001110010";
                when x"E8" => data <= "0000000001";
                when x"E9" => data <= "1100111011";
                when x"EA" => data <= "1111011010";
                when x"EB" => data <= "1111011010";
                when x"EC" => data <= "1111101111";
                when x"ED" => data <= "0000000001";
                when x"EE" => data <= "1111101111";
                when x"EF" => data <= "0010001010";
                when x"F0" => data <= "1111011010";
                when x"F1" => data <= "1000101101";
                when x"F2" => data <= "1111101111";
                when x"F3" => data <= "0110011100";
                when x"F4" => data <= "1111011010";
                when x"F5" => data <= "0010001010";
                when x"F6" => data <= "0000000001";
                when x"F7" => data <= "1111011010";
                when x"F8" => data <= "1011111001";
                when x"F9" => data <= "1111011010";
                when x"FA" => data <= "0000000001";
                when x"FB" => data <= "0110101001";
                when x"FC" => data <= "0101111101";
                when x"FD" => data <= "1111011010";
                when x"FE" => data <= "1111011010";
                when x"FF" => data <= "0100100010";
                when x"100" => data <= "0010111111";
                when x"101" => data <= "1001000111";
                when x"102" => data <= "1111011010";
                when x"103" => data <= "1111011010";
                when x"104" => data <= "1000011000";
                when x"105" => data <= "0110011100";
                when x"106" => data <= "1111011010";
                when x"107" => data <= "0100010111";
                when x"108" => data <= "1000101101";
                when x"109" => data <= "0000000001";
                when x"10A" => data <= "0000000001";
                when x"10B" => data <= "0110101001";
                when x"10C" => data <= "1100111011";
                when x"10D" => data <= "1100111011";
                when x"10E" => data <= "0010001010";
                when x"10F" => data <= "1111101111";
                when x"110" => data <= "1000101101";
                when x"111" => data <= "1100001110";
                when x"112" => data <= "1000101101";
                when x"113" => data <= "1111011010";
                when x"114" => data <= "1111011010";
                when x"115" => data <= "1111011010";
                when x"116" => data <= "0000000001";
                when x"117" => data <= "0111111101";
                when x"118" => data <= "0010000001";
                when x"119" => data <= "0000001010";
                when x"11A" => data <= "0111111101";
                when x"11B" => data <= "1101011010";
                when x"11C" => data <= "1101011010";
                when x"11D" => data <= "0110100010";
                when x"11E" => data <= "1010101101";
                when x"11F" => data <= "1110111011";
                when x"120" => data <= "0000111111";
                when x"121" => data <= "1101011010";
                when x"122" => data <= "0111001000";
                when x"123" => data <= "1010101101";
                when x"124" => data <= "0000111111";
                when x"125" => data <= "1010101101";
                when x"126" => data <= "1010101101";
                when x"127" => data <= "1110111011";
                when x"128" => data <= "1010011000";
                when x"129" => data <= "0111001000";
                when x"12A" => data <= "0100101001";
                when x"12B" => data <= "0111001000";
                when x"12C" => data <= "1110001110";
                when x"12D" => data <= "1100110000";
                when x"12E" => data <= "0100101001";
                when x"12F" => data <= "0111001000";
                when x"130" => data <= "0000001010";
                when x"131" => data <= "1010011000";
                when x"132" => data <= "0111111101";
                when x"133" => data <= "1101011010";
                when x"134" => data <= "0011101011";
                when x"135" => data <= "1010101101";
                when x"136" => data <= "0111111101";
                when x"137" => data <= "1110111011";
                when x"138" => data <= "1010101101";
                when x"139" => data <= "0100101001";
                when x"13A" => data <= "1110111011";
                when x"13B" => data <= "1110111011";
                when x"13C" => data <= "0001010101";
                when x"13D" => data <= "1111111110";
                when x"13E" => data <= "1011101000";
                when x"13F" => data <= "1111111110";
                when x"140" => data <= "0000010000";
                when x"141" => data <= "0000100101";
                when x"142" => data <= "1111111110";
                when x"143" => data <= "0001001111";
                when x"144" => data <= "0111100111";
                when x"145" => data <= "0111100111";
                when x"146" => data <= "0100000110";
                when x"147" => data <= "0100110011";
                when x"148" => data <= "0000100101";
                when x"149" => data <= "1000001001";
                when x"14A" => data <= "1000001001";
                when x"14B" => data <= "0000100101";
                when x"14C" => data <= "0100000110";
                when x"14D" => data <= "0000100101";
                when x"14E" => data <= "1010000010";
                when x"14F" => data <= "0111100111";
                when x"150" => data <= "0000010000";
                when x"151" => data <= "0111010010";
                when x"152" => data <= "0100000110";
                when x"153" => data <= "1111111110";
                when x"154" => data <= "1111111110";
                when x"155" => data <= "0000100101";
                when x"156" => data <= "0000100101";
                when x"157" => data <= "0111010010";
                when x"158" => data <= "1111111110";
                when x"159" => data <= "0110001101";
                when x"15A" => data <= "1011101000";
                when x"15B" => data <= "0000010000";
                when x"15C" => data <= "0000100101";
                when x"15D" => data <= "0000100101";
                when x"15E" => data <= "1111111110";
                when x"15F" => data <= "0001111010";
                when x"160" => data <= "1111111110";
                when x"161" => data <= "0100000110";
                when x"162" => data <= "1111111110";
                when x"163" => data <= "0000100101";
                when x"164" => data <= "0111100111";
                when x"165" => data <= "0111100111";
                when x"166" => data <= "1111111110";
                when x"167" => data <= "1111111110";
                when x"168" => data <= "0000100101";
                when x"169" => data <= "0000100101";
                when x"16A" => data <= "0100000110";
                when x"16B" => data <= "1000111100";
                when x"16C" => data <= "0011000100";
                when x"16D" => data <= "1000001001";
                when x"16E" => data <= "1111111110";
                when x"16F" => data <= "1111111110";
                when x"170" => data <= "0000010000";
                when x"171" => data <= "0000100101";
                when x"172" => data <= "0111010010";
                when x"173" => data <= "0000100101";
                when x"174" => data <= "1111111110";
                when x"175" => data <= "1000001001";
                when x"176" => data <= "0000100101";
                when x"177" => data <= "1111111110";
                when x"178" => data <= "1111111110";
                when x"179" => data <= "0000100101";
                when x"17A" => data <= "0011000100";
                when x"17B" => data <= "0000010000";
                when x"17C" => data <= "0100110011";
                when x"17D" => data <= "1111111110";
                when x"17E" => data <= "0000100101";
                when x"17F" => data <= "0000010000";
                when x"180" => data <= "0110011010";
                when x"181" => data <= "0100100100";
                when x"182" => data <= "1011111111";
                when x"183" => data <= "1011111111";
                when x"184" => data <= "1011111111";
                when x"185" => data <= "1011111111";
                when x"186" => data <= "1011111111";
                when x"187" => data <= "0110101111";
                when x"188" => data <= "0110101111";
                when x"189" => data <= "1011111111";
                when x"18A" => data <= "1011111111";
                when x"18B" => data <= "1011111111";
                when x"18C" => data <= "0001011000";
                when x"18D" => data <= "1011111111";
                when x"18E" => data <= "1011111111";
                when x"18F" => data <= "1011111111";
                when x"190" => data <= "1011111111";
                when x"191" => data <= "0001101101";
                when x"192" => data <= "1001000001";
                when x"193" => data <= "1011111111";
                when x"194" => data <= "1011111111";
                when x"195" => data <= "0001101101";
                when x"196" => data <= "1011111111";
                when x"197" => data <= "1011111111";
                when x"198" => data <= "1011111111";
                when x"199" => data <= "1011111111";
                when x"19A" => data <= "1011111111";
                when x"19B" => data <= "1011111111";
                when x"19C" => data <= "1011111111";
                when x"19D" => data <= "1011111111";
                when x"19E" => data <= "1011111111";
                when x"19F" => data <= "1011111111";
                when x"1A0" => data <= "0010001100";
                when x"1A1" => data <= "1011111111";
                when x"1A2" => data <= "1011111111";
                when x"1A3" => data <= "1011111111";
                when x"1A4" => data <= "1011111111";
                when x"1A5" => data <= "1011111111";
                when x"1A6" => data <= "1011111111";
                when x"1A7" => data <= "1011111111";
                when x"1A8" => data <= "1011111111";
                when x"1A9" => data <= "0110101111";
                when x"1AA" => data <= "1011111111";
                when x"1AB" => data <= "1011111111";
                when x"1AC" => data <= "1011111111";
                when x"1AD" => data <= "1011111111";
                when x"1AE" => data <= "1011111111";
                when x"1AF" => data <= "1011111111";
                when x"1B0" => data <= "1100001000";
                when x"1B1" => data <= "1101010111";
                when x"1B2" => data <= "1011111111";
                when x"1B3" => data <= "0001011000";
                when x"1B4" => data <= "1011111111";
                when x"1B5" => data <= "1010100000";
                when x"1B6" => data <= "1110110110";
                when x"1B7" => data <= "0110011010";
                when x"1B8" => data <= "0010001100";
                when x"1B9" => data <= "0101111011";
                when x"1BA" => data <= "1011111111";
                when x"1BB" => data <= "1011111111";
                when x"1BC" => data <= "1011111111";
                when x"1BD" => data <= "1011111111";
                when x"1BE" => data <= "1011111111";
                when x"1BF" => data <= "1011111111";
                when x"1C0" => data <= "1011111111";
                when x"1C1" => data <= "1011111111";
                when x"1C2" => data <= "1011111111";
                when x"1C3" => data <= "1011111111";
                when x"1C4" => data <= "0100100100";
                when x"1C5" => data <= "0001101101";
                when x"1C6" => data <= "1011111111";
                when x"1C7" => data <= "1011001010";
                when x"1C8" => data <= "1011111111";
                when x"1C9" => data <= "1011111111";
                when x"1CA" => data <= "1101010111";
                when x"1CB" => data <= "1011111111";
                when x"1CC" => data <= "0110101111";
                when x"1CD" => data <= "0000000111";
                when x"1CE" => data <= "1011111111";
                when x"1CF" => data <= "1011111111";
                when x"1D0" => data <= "1011111111";
                when x"1D1" => data <= "0110101111";
                when x"1D2" => data <= "1011111111";
                when x"1D3" => data <= "1011111111";
                when x"1D4" => data <= "1011111111";
                when x"1D5" => data <= "1011111111";
                when x"1D6" => data <= "1011111111";
                when x"1D7" => data <= "1011111111";
                when x"1D8" => data <= "1011111111";
                when x"1D9" => data <= "1011111111";
                when x"1DA" => data <= "1011111111";
                when x"1DB" => data <= "0101111011";
                when x"1DC" => data <= "1011111111";
                when x"1DD" => data <= "1011111111";
                when x"1DE" => data <= "0110011010";
                when x"1DF" => data <= "0110101111";
                when x"1E0" => data <= "1011111111";
                when x"1E1" => data <= "1011111111";
                when x"1E2" => data <= "1011111111";
                when x"1E3" => data <= "1011111111";
                when x"1E4" => data <= "0110101111";
                when x"1E5" => data <= "1011111111";
                when x"1E6" => data <= "1011111111";
                when x"1E7" => data <= "1100111101";
                when x"1E8" => data <= "1011111111";
                when x"1E9" => data <= "1011111111";
                when x"1EA" => data <= "1011111111";
                when x"1EB" => data <= "1011111111";
                when x"1EC" => data <= "1011111111";
                when x"1ED" => data <= "1011111111";
                when x"1EE" => data <= "1011111111";
                when x"1EF" => data <= "1010100000";
                when x"1F0" => data <= "1011111111";
                when x"1F1" => data <= "1011111111";
                when x"1F2" => data <= "1011111111";
                when x"1F3" => data <= "1011111111";
                when x"1F4" => data <= "1011111111";
                when x"1F5" => data <= "0110101111";
                when x"1F6" => data <= "1011111111";
                when x"1F7" => data <= "1011111111";
                when x"1F8" => data <= "1011111111";
                when x"1F9" => data <= "0110101111";
                when x"1FA" => data <= "1101010111";
                when x"1FB" => data <= "1011111111";
                when x"1FC" => data <= "1011111111";
                when x"1FD" => data <= "1101111000";
                when x"1FE" => data <= "0110000000";
                when x"1FF" => data <= "0100001011";
                when x"200" => data <= "0110000000";
                when x"201" => data <= "0110000000";
                when x"202" => data <= "1000000100";
                when x"203" => data <= "0111011111";
                when x"204" => data <= "1000110001";
                when x"205" => data <= "1111110011";
                when x"206" => data <= "0001000010";
                when x"207" => data <= "0110000000";
                when x"208" => data <= "0000101000";
                when x"209" => data <= "0000101000";
                when x"20A" => data <= "0110000000";
                when x"20B" => data <= "0110000000";
                when x"20C" => data <= "1100100111";
                when x"20D" => data <= "0111011111";
                when x"20E" => data <= "1000000100";
                when x"20F" => data <= "0111011111";
                when x"210" => data <= "1000000100";
                when x"211" => data <= "0000101000";
                when x"212" => data <= "0101010100";
                when x"213" => data <= "1000000100";
                when x"214" => data <= "1011010000";
                when x"215" => data <= "1000000100";
                when x"216" => data <= "0111011111";
                when x"217" => data <= "1000110001";
                when x"218" => data <= "1001011011";
                when x"219" => data <= "0001000010";
                when x"21A" => data <= "0010100011";
                when x"21B" => data <= "1011010000";
                when x"21C" => data <= "0111011111";
                when x"21D" => data <= "0000101000";
                when x"21E" => data <= "1000000100";
                when x"21F" => data <= "0110000000";
                when x"220" => data <= "1000000100";
                when x"221" => data <= "1000000100";
                when x"222" => data <= "0110000000";
                when x"223" => data <= "1111110011";
                when x"224" => data <= "0000101000";
                when x"225" => data <= "0001000010";
                when x"226" => data <= "1000000100";
                when x"227" => data <= "1000000100";
                when x"228" => data <= "0000101000";
                when x"229" => data <= "0111011111";
                when x"22A" => data <= "0101010100";
                when x"22B" => data <= "0111011111";
                when x"22C" => data <= "0100001011";
                when x"22D" => data <= "1011010000";
                when x"22E" => data <= "0110000000";
                when x"22F" => data <= "1001011011";
                when x"230" => data <= "0110000000";
                when x"231" => data <= "0110000000";
                when x"232" => data <= "1000000100";
                when x"233" => data <= "0111011111";
                when x"234" => data <= "0110000000";
                when x"235" => data <= "0111011111";
                when x"236" => data <= "0110000000";
                when x"237" => data <= "1000000100";
                when x"238" => data <= "0001000010";
                when x"239" => data <= "0111011111";
                when x"23A" => data <= "1000000100";
                when x"23B" => data <= "1000000100";
                when x"23C" => data <= "1000000100";
                when x"23D" => data <= "0111011111";
                when x"23E" => data <= "0000101000";
                when x"23F" => data <= "1000000100";
                when x"240" => data <= "0000101000";
                when x"241" => data <= "1000000100";
                when x"242" => data <= "1111110110";
                when x"243" => data <= "1010111111";
                when x"244" => data <= "0111011010";
                when x"245" => data <= "0111101111";
                when x"246" => data <= "1010001010";
                when x"247" => data <= "1010111111";
                when x"248" => data <= "0000101101";
                when x"249" => data <= "0111011010";
                when x"24A" => data <= "1010111111";
                when x"24B" => data <= "0000101101";
                when x"24C" => data <= "1010111111";
                when x"24D" => data <= "0111011010";
                when x"24E" => data <= "0100111011";
                when x"24F" => data <= "0111101111";
                when x"250" => data <= "0000011000";
                when x"251" => data <= "1000110100";
                when x"252" => data <= "0000011000";
                when x"253" => data <= "1010001010";
                when x"254" => data <= "0000101101";
                when x"255" => data <= "0000101101";
                when x"256" => data <= "0111101111";
                when x"257" => data <= "0000101101";
                when x"258" => data <= "1111110110";
                when x"259" => data <= "1000000001";
                when x"25A" => data <= "1010111111";
                when x"25B" => data <= "0000101101";
                when x"25C" => data <= "1010111111";
                when x"25D" => data <= "1101111101";
                when x"25E" => data <= "0000101101";
                when x"25F" => data <= "1010111111";
                when x"260" => data <= "0000101101";
                when x"261" => data <= "0111101111";
                when x"262" => data <= "0000011000";
                when x"263" => data <= "0111011010";
                when x"264" => data <= "1000000001";
                when x"265" => data <= "1101111101";
                when x"266" => data <= "1010111111";
                when x"267" => data <= "1010111111";
                when x"268" => data <= "0111101111";
                when x"269" => data <= "1110011100";
                when x"26A" => data <= "1101111101";
                when x"26B" => data <= "0000101101";
                when x"26C" => data <= "0111101111";
                when x"26D" => data <= "0111101111";
                when x"26E" => data <= "0111011010";
                when x"26F" => data <= "0111101111";
                when x"270" => data <= "0100111011";
                when x"271" => data <= "1101111101";
                when x"272" => data <= "1101111101";
                when x"273" => data <= "1010111111";
                when x"274" => data <= "1010111111";
                when x"275" => data <= "1101111101";
                when x"276" => data <= "0111101111";
                when x"277" => data <= "0111011010";
                when x"278" => data <= "0000011000";
                when x"279" => data <= "0001000111";
                when x"27A" => data <= "0111101111";
                when x"27B" => data <= "0000101101";
                when x"27C" => data <= "0111101111";
                when x"27D" => data <= "1010111111";
                when x"27E" => data <= "0111101111";
                when x"27F" => data <= "1000000001";
                when x"280" => data <= "0100111011";
                when x"281" => data <= "0111101111";
                when x"282" => data <= "1010111111";
                when x"283" => data <= "0111101111";
                when x"284" => data <= "1000110100";
                when x"285" => data <= "1000000001";
                when x"286" => data <= "1101111101";
                when x"287" => data <= "1010001010";
                when x"288" => data <= "1101010010";
                when x"289" => data <= "1001110001";
                when x"28A" => data <= "0000000010";
                when x"28B" => data <= "0000000010";
                when x"28C" => data <= "0000000010";
                when x"28D" => data <= "1110000110";
                when x"28E" => data <= "0000000010";
                when x"28F" => data <= "0000000010";
                when x"290" => data <= "1001000100";
                when x"291" => data <= "0000000010";
                when x"292" => data <= "0000000010";
                when x"293" => data <= "0111110101";
                when x"294" => data <= "1011111010";
                when x"295" => data <= "1011111010";
                when x"296" => data <= "1001110001";
                when x"297" => data <= "1101010010";
                when x"298" => data <= "0111000000";
                when x"299" => data <= "1101010010";
                when x"29A" => data <= "1011111010";
                when x"29B" => data <= "0100010100";
                when x"29C" => data <= "0110101010";
                when x"29D" => data <= "1010100101";
                when x"29E" => data <= "1010100101";
                when x"29F" => data <= "0000000010";
                when x"2A0" => data <= "0100010100";
                when x"2A1" => data <= "1011111010";
                when x"2A2" => data <= "0111110101";
                when x"2A3" => data <= "0111000000";
                when x"2A4" => data <= "0000000010";
                when x"2A5" => data <= "0111000000";
                when x"2A6" => data <= "0111000000";
                when x"2A7" => data <= "1100001101";
                when x"2A8" => data <= "0000000010";
                when x"2A9" => data <= "1010100101";
                when x"2AA" => data <= "0110011111";
                when x"2AB" => data <= "0000000010";
                when x"2AC" => data <= "0000000010";
                when x"2AD" => data <= "0011010110";
                when x"2AE" => data <= "0100010100";
                when x"2AF" => data <= "1110000110";
                when x"2B0" => data <= "0000000010";
                when x"2B1" => data <= "1001110001";
                when x"2B2" => data <= "0110101010";
                when x"2B3" => data <= "0110011111";
                when x"2B4" => data <= "1001000100";
                when x"2B5" => data <= "1111011001";
                when x"2B6" => data <= "1011111010";
                when x"2B7" => data <= "1111111011";
                when x"2B8" => data <= "1111111011";
                when x"2B9" => data <= "0110001000";
                when x"2BA" => data <= "1111111011";
                when x"2BB" => data <= "1111111011";
                when x"2BC" => data <= "1111111011";
                when x"2BD" => data <= "0111010111";
                when x"2BE" => data <= "1000111001";
                when x"2BF" => data <= "0000100000";
                when x"2C0" => data <= "1000111001";
                when x"2C1" => data <= "0000100000";
                when x"2C2" => data <= "1011011000";
                when x"2C3" => data <= "0110001000";
                when x"2C4" => data <= "0000100000";
                when x"2C5" => data <= "1000111001";
                when x"2C6" => data <= "1011011000";
                when x"2C7" => data <= "0000010101";
                when x"2C8" => data <= "1111111011";
                when x"2C9" => data <= "0000100000";
                when x"2CA" => data <= "0110001000";
                when x"2CB" => data <= "1111111011";
                when x"2CC" => data <= "0111010111";
                when x"2CD" => data <= "1111111011";
                when x"2CE" => data <= "1111111011";
                when x"2CF" => data <= "1011101101";
                when x"2D0" => data <= "0110001000";
                when x"2D1" => data <= "0100000011";
                when x"2D2" => data <= "1011011000";
                when x"2D3" => data <= "0100000011";
                when x"2D4" => data <= "1111111011";
                when x"2D5" => data <= "0000100000";
                when x"2D6" => data <= "0010101011";
                when x"2D7" => data <= "1111111011";
                when x"2D8" => data <= "0000100000";
                when x"2D9" => data <= "1111111011";
                when x"2DA" => data <= "0000100000";
                when x"2DB" => data <= "0001111111";
                when x"2DC" => data <= "0000100000";
                when x"2DD" => data <= "0000010101";
                when x"2DE" => data <= "1111111011";
                when x"2DF" => data <= "1111111011";
                when x"2E0" => data <= "1111111011";
                when x"2E1" => data <= "1111111011";
                when x"2E2" => data <= "1111111011";
                when x"2E3" => data <= "0000100000";
                when x"2E4" => data <= "0000100000";
                when x"2E5" => data <= "0000100000";
                when x"2E6" => data <= "0000100000";
                when x"2E7" => data <= "0110001000";
                when x"2E8" => data <= "0000100000";
                when x"2E9" => data <= "0110001000";
                when x"2EA" => data <= "0001001010";
                when x"2EB" => data <= "1111111011";
                when x"2EC" => data <= "0000100000";
                when x"2ED" => data <= "0111010111";
                when x"2EE" => data <= "1111111011";
                when x"2EF" => data <= "1111111011";
                when x"2F0" => data <= "1011101101";
                when x"2F1" => data <= "1111111011";
                when x"2F2" => data <= "0111100010";
                when x"2F3" => data <= "0000100000";
                when x"2F4" => data <= "1111111011";
                when x"2F5" => data <= "0000100000";
                when x"2F6" => data <= "1111111011";
                when x"2F7" => data <= "1111111011";
                when x"2F8" => data <= "1111111011";
                when x"2F9" => data <= "1111111011";
                when x"2FA" => data <= "0000100000";
                when x"2FB" => data <= "0010101011";
                when x"2FC" => data <= "1111111011";
                when x"2FD" => data <= "0000100000";
                when x"2FE" => data <= "1111111011";
                when x"2FF" => data <= "1111111011";
                when x"300" => data <= "0000100000";
                when x"301" => data <= "1100011010";
                when x"302" => data <= "1111111011";
                when x"303" => data <= "0000100000";
                when x"304" => data <= "1111111011";
                when x"305" => data <= "1111111011";
                when x"306" => data <= "1111111011";
                when x"307" => data <= "0000100000";
                when x"308" => data <= "0000100000";
                when x"309" => data <= "1011011000";
                when x"30A" => data <= "1111111011";
                when x"30B" => data <= "1100101111";
                when x"30C" => data <= "1111111011";
                when x"30D" => data <= "1000111001";
                when x"30E" => data <= "1111111011";
                when x"30F" => data <= "1111111011";
                when x"310" => data <= "1111111011";
                when x"311" => data <= "1011000010";
                when x"312" => data <= "0001010000";
                when x"313" => data <= "1000010110";
                when x"314" => data <= "1111010100";
                when x"315" => data <= "1011110111";
                when x"316" => data <= "1111010100";
                when x"317" => data <= "0101000110";
                when x"318" => data <= "1100000000";
                when x"319" => data <= "0101110011";
                when x"31A" => data <= "1011110111";
                when x"31B" => data <= "1001001001";
                when x"31C" => data <= "1011110111";
                when x"31D" => data <= "1110001011";
                when x"31E" => data <= "1010101000";
                when x"31F" => data <= "1000010110";
                when x"320" => data <= "1000100011";
                when x"321" => data <= "0001010000";
                when x"322" => data <= "0001010000";
                when x"323" => data <= "0001010000";
                when x"324" => data <= "1010101000";
                when x"325" => data <= "0001010000";
                when x"326" => data <= "0001010000";
                when x"327" => data <= "1100000000";
                when x"328" => data <= "0110100111";
                when x"329" => data <= "1101011111";
                when x"32A" => data <= "1101011111";
                when x"32B" => data <= "0010000100";
                when x"32C" => data <= "0110100111";
                when x"32D" => data <= "1100000000";
                when x"32E" => data <= "0001100101";
                when x"32F" => data <= "1010101000";
                when x"330" => data <= "1011110111";
                when x"331" => data <= "0001010000";
                when x"332" => data <= "0110100111";
                when x"333" => data <= "1011110111";
                when x"334" => data <= "0010000100";
                when x"335" => data <= "1110111110";
                when x"336" => data <= "0110100111";
                when x"337" => data <= "1010101000";
                when x"338" => data <= "1010101000";
                when x"339" => data <= "1100000000";
                when x"33A" => data <= "1011110111";
                when x"33B" => data <= "1101011111";
                when x"33C" => data <= "1011110111";
                when x"33D" => data <= "1100110101";
                when x"33E" => data <= "1101011111";
                when x"33F" => data <= "0101000110";
                when x"340" => data <= "0010000100";
                when x"341" => data <= "1000100011";
                when x"342" => data <= "1011110111";
                when x"343" => data <= "1001000010";
                when x"344" => data <= "0000000100";
                when x"345" => data <= "0000000100";
                when x"346" => data <= "1111011111";
                when x"347" => data <= "0000000100";
                when x"348" => data <= "1001000010";
                when x"349" => data <= "1111011111";
                when x"34A" => data <= "1111011111";
                when x"34B" => data <= "1001110111";
                when x"34C" => data <= "1111011111";
                when x"34D" => data <= "0111000110";
                when x"34E" => data <= "1111011111";
                when x"34F" => data <= "0000000100";
                when x"350" => data <= "0000000100";
                when x"351" => data <= "0111000110";
                when x"352" => data <= "1001110111";
                when x"353" => data <= "0000000100";
                when x"354" => data <= "0000000100";
                when x"355" => data <= "0000000100";
                when x"356" => data <= "1000101000";
                when x"357" => data <= "0000000100";
                when x"358" => data <= "0000000100";
                when x"359" => data <= "1111011111";
                when x"35A" => data <= "0000000100";
                when x"35B" => data <= "1001000010";
                when x"35C" => data <= "1111011111";
                when x"35D" => data <= "0000000100";
                when x"35E" => data <= "0000000100";
                when x"35F" => data <= "0000000100";
                when x"360" => data <= "1000101000";
                when x"361" => data <= "0000000100";
                when x"362" => data <= "0000000100";
                when x"363" => data <= "1110110101";
                when x"364" => data <= "1001000010";
                when x"365" => data <= "1110000000";
                when x"366" => data <= "0000000100";
                when x"367" => data <= "0000000100";
                when x"368" => data <= "0000000100";
                when x"369" => data <= "1111011111";
                when x"36A" => data <= "1111011111";
                when x"36B" => data <= "1111011111";
                when x"36C" => data <= "0000000100";
                when x"36D" => data <= "0111000110";
                when x"36E" => data <= "0100010010";
                when x"36F" => data <= "1001000010";
                when x"370" => data <= "0000000100";
                when x"371" => data <= "1111101010";
                when x"372" => data <= "0010111010";
                when x"373" => data <= "1001110111";
                when x"374" => data <= "1110000000";
                when x"375" => data <= "1101010100";
                when x"376" => data <= "0000000100";
                when x"377" => data <= "0000000100";
                when x"378" => data <= "0100010010";
                when x"379" => data <= "1111011111";
                when x"37A" => data <= "0000000100";
                when x"37B" => data <= "1111011111";
                when x"37C" => data <= "0000000100";
                when x"37D" => data <= "0000000100";
                when x"37E" => data <= "1111011111";
                when x"37F" => data <= "0000000100";
                when x"380" => data <= "1000101000";
                when x"381" => data <= "0000000100";
                when x"382" => data <= "0011100101";
                when x"383" => data <= "0000000100";
                when x"384" => data <= "1001000010";
                when x"385" => data <= "0000000100";
                when x"386" => data <= "1111011111";
                when x"387" => data <= "0000000100";
                when x"388" => data <= "0100100111";
                when x"389" => data <= "0000000100";
                when x"38A" => data <= "0000000100";
                when x"38B" => data <= "1001110111";
                when x"38C" => data <= "0100010010";
                when x"38D" => data <= "0000000100";
                when x"38E" => data <= "1001110111";
                when x"38F" => data <= "1110000000";
                when x"390" => data <= "1001110111";
                when x"391" => data <= "1111011111";
                when x"392" => data <= "0000000100";
                when x"393" => data <= "1110000000";
                when x"394" => data <= "0000000100";
                when x"395" => data <= "1001110111";
                when x"396" => data <= "0000000100";
                when x"397" => data <= "1000101000";
                when x"398" => data <= "1111011111";
                when x"399" => data <= "1000011101";
                when x"39A" => data <= "1001000010";
                when x"39B" => data <= "0000000100";
                when x"39C" => data <= "0000000100";
                when x"39D" => data <= "0000000100";
                when x"39E" => data <= "0110101100";
                when x"39F" => data <= "0011111111";
                when x"3A0" => data <= "1001011000";
                when x"3A1" => data <= "0011111111";
                when x"3A2" => data <= "0100001000";
                when x"3A3" => data <= "0100001000";
                when x"3A4" => data <= "0011001010";
                when x"3A5" => data <= "0100111101";
                when x"3A6" => data <= "0000101011";
                when x"3A7" => data <= "1001011000";
                when x"3A8" => data <= "0011111111";
                when x"3A9" => data <= "1110101111";
                when x"3AA" => data <= "0100001000";
                when x"3AB" => data <= "1110011010";
                when x"3AC" => data <= "0100001000";
                when x"3AD" => data <= "0100001000";
                when x"3AE" => data <= "1001011000";
                when x"3AF" => data <= "1110011010";
                when x"3B0" => data <= "1001011000";
                when x"3B1" => data <= "0101100010";
                when x"3B2" => data <= "1110101111";
                when x"3B3" => data <= "0100001000";
                when x"3B4" => data <= "1010111001";
                when x"3B5" => data <= "1001011000";
                when x"3B6" => data <= "0010100000";
                when x"3B7" => data <= "1110101111";
                when x"3B8" => data <= "1110101111";
                when x"3B9" => data <= "1101111011";
                when x"3BA" => data <= "1101111011";
                when x"3BB" => data <= "0100111101";
                when x"3BC" => data <= "0101010111";
                when x"3BD" => data <= "0011111111";
                when x"3BE" => data <= "1001011000";
                when x"3BF" => data <= "1110101111";
                when x"3C0" => data <= "0011111111";
                when x"3C1" => data <= "1111110000";
                when x"3C2" => data <= "0011111111";
                when x"3C3" => data <= "0100111101";
                when x"3C4" => data <= "1101111011";
                when x"3C5" => data <= "0100001000";
                when x"3C6" => data <= "1101111011";
                when x"3C7" => data <= "0100001000";
                when x"3C8" => data <= "0011001010";
                when x"3C9" => data <= "1110101111";
                when x"3CA" => data <= "0011111111";
                when x"3CB" => data <= "0101010111";
                when x"3CC" => data <= "0100001000";
                when x"3CD" => data <= "0011001010";
                when x"3CE" => data <= "0100001000";
                when x"3CF" => data <= "1101111011";
                when x"3D0" => data <= "1011010011";
                when x"3D1" => data <= "0011111111";
                when x"3D2" => data <= "0100001000";
                when x"3D3" => data <= "0001000001";
                when x"3D4" => data <= "0011001010";
                when x"3D5" => data <= "0011001010";
                when x"3D6" => data <= "1000000111";
                when x"3D7" => data <= "0100111101";
                when x"3D8" => data <= "1110101111";
                when x"3D9" => data <= "0101000000";
                when x"3DA" => data <= "1000010000";
                when x"3DB" => data <= "0111111110";
                when x"3DC" => data <= "1000010000";
                when x"3DD" => data <= "1111010010";
                when x"3DE" => data <= "0101000000";
                when x"3DF" => data <= "1110111000";
                when x"3E0" => data <= "1111010010";
                when x"3E1" => data <= "1000010000";
                when x"3E2" => data <= "1100000110";
                when x"3E3" => data <= "0101000000";
                when x"3E4" => data <= "1110111000";
                when x"3E5" => data <= "1000010000";
                when x"3E6" => data <= "0101110101";
                when x"3E7" => data <= "1110111000";
                when x"3E8" => data <= "0111111110";
                when x"3E9" => data <= "1000100101";
                when x"3EA" => data <= "1011110001";
                when x"3EB" => data <= "0010000010";
                when x"3EC" => data <= "1101011001";
                when x"3ED" => data <= "0101000000";
                when x"3EE" => data <= "1000010000";
                when x"3EF" => data <= "0101110101";
                when x"3F0" => data <= "0101000000";
                when x"3F1" => data <= "0000001001";
                when x"3F2" => data <= "1000010000";
                when x"3F3" => data <= "1000010000";
                when x"3F4" => data <= "0101110101";
                when x"3F5" => data <= "0101000000";
                when x"3F6" => data <= "1111010010";
                when x"3F7" => data <= "1001111010";
                when x"3F8" => data <= "1110111000";
                when x"3F9" => data <= "1000010000";
                when x"3FA" => data <= "1111100111";
                when x"3FB" => data <= "1111010010";
                when x"3FC" => data <= "1000100101";
                when x"3FD" => data <= "0101000000";
                when x"3FE" => data <= "1000010000";
                when x"3FF" => data <= "1010101110";
                when x"400" => data <= "1111010010";
                when x"401" => data <= "1111010010";
                when x"402" => data <= "0001010110";
                when x"403" => data <= "0101000000";
                when x"404" => data <= "0010000010";
                when x"405" => data <= "0111001011";
                when x"406" => data <= "1000010000";
                when x"407" => data <= "0101110101";
                when x"408" => data <= "0101110101";
                when x"409" => data <= "0101110101";
                when x"40A" => data <= "1110111000";
                when x"40B" => data <= "0111001011";
                when x"40C" => data <= "1000010000";
                when x"40D" => data <= "0101000000";
                when x"40E" => data <= "0010000010";
                when x"40F" => data <= "0101110101";
                when x"410" => data <= "0101110101";
                when x"411" => data <= "0010000010";
                when x"412" => data <= "1010101110";
                when x"413" => data <= "1000100101";
                when x"414" => data <= "0101110101";
                when x"415" => data <= "0101110101";
                when x"416" => data <= "0101000000";
                when x"417" => data <= "0001010110";
                when x"418" => data <= "1000010000";
                when x"419" => data <= "1000100101";
                when x"41A" => data <= "1111111101";
                when x"41B" => data <= "0011110010";
                when x"41C" => data <= "0000010011";
                when x"41D" => data <= "1111001000";
                when x"41E" => data <= "0101011010";
                when x"41F" => data <= "1000111111";
                when x"420" => data <= "1011011110";
                when x"421" => data <= "1111111101";
                when x"422" => data <= "1111111101";
                when x"423" => data <= "0100000101";
                when x"424" => data <= "1110010111";
                when x"425" => data <= "1000111111";
                when x"426" => data <= "0101101111";
                when x"427" => data <= "1000001010";
                when x"428" => data <= "1011011110";
                when x"429" => data <= "0100000101";
                when x"42A" => data <= "1000001010";
                when x"42B" => data <= "1001010101";
                when x"42C" => data <= "1111001000";
                when x"42D" => data <= "1111111101";
                when x"42E" => data <= "1111001000";
                when x"42F" => data <= "1111111101";
                when x"430" => data <= "1011101011";
                when x"431" => data <= "0010011000";
                when x"432" => data <= "1111111101";
                when x"433" => data <= "1111111101";
                when x"434" => data <= "1011011110";
                when x"435" => data <= "0111010001";
                when x"436" => data <= "0100000101";
                when x"437" => data <= "1111111101";
                when x"438" => data <= "0001001100";
                when x"439" => data <= "1111111101";
                when x"43A" => data <= "0100000101";
                when x"43B" => data <= "1111111101";
                when x"43C" => data <= "1110010111";
                when x"43D" => data <= "1111111101";
                when x"43E" => data <= "1111111101";
                when x"43F" => data <= "1000111111";
                when x"440" => data <= "1111111101";
                when x"441" => data <= "1001010101";
                when x"442" => data <= "0101101111";
                when x"443" => data <= "1000001010";
                when x"444" => data <= "1000111111";
                when x"445" => data <= "1111111101";
                when x"446" => data <= "0100000101";
                when x"447" => data <= "0010101101";
                when x"448" => data <= "0100000101";
                when x"449" => data <= "1001100000";
                when x"44A" => data <= "1111111101";
                when x"44B" => data <= "1111111101";
                when x"44C" => data <= "1100111111";
                when x"44D" => data <= "1010100010";
                when x"44E" => data <= "1010010111";
                when x"44F" => data <= "1111011110";
                when x"450" => data <= "1100111111";
                when x"451" => data <= "1011111101";
                when x"452" => data <= "0010111011";
                when x"453" => data <= "1111011110";
                when x"454" => data <= "0110101101";
                when x"455" => data <= "0111000111";
                when x"456" => data <= "1100111111";
                when x"457" => data <= "0000000101";
                when x"458" => data <= "1011111101";
                when x"459" => data <= "0110101101";
                when x"45A" => data <= "1100111111";
                when x"45B" => data <= "0000000101";
                when x"45C" => data <= "1000011100";
                when x"45D" => data <= "1011111101";
                when x"45E" => data <= "1011111101";
                when x"45F" => data <= "0110101101";
                when x"460" => data <= "1110110100";
                when x"461" => data <= "0110101101";
                when x"462" => data <= "0000000101";
                when x"463" => data <= "0000000101";
                when x"464" => data <= "1011111101";
                when x"465" => data <= "1000101001";
                when x"466" => data <= "1111011110";
                when x"467" => data <= "1011111101";
                when x"468" => data <= "1100111111";
                when x"469" => data <= "0000000101";
                when x"46A" => data <= "1100111111";
                when x"46B" => data <= "0000000101";
                when x"46C" => data <= "0000000101";
                when x"46D" => data <= "0110101101";
                when x"46E" => data <= "1011001000";
                when x"46F" => data <= "0110011000";
                when x"470" => data <= "1100111111";
                when x"471" => data <= "1100111111";
                when x"472" => data <= "1011001000";
                when x"473" => data <= "0110101101";
                when x"474" => data <= "1010100010";
                when x"475" => data <= "0000000101";
                when x"476" => data <= "1000101001";
                when x"477" => data <= "1100111111";
                when x"478" => data <= "1111011110";
                when x"479" => data <= "0000000101";
                when x"47A" => data <= "1111011110";
                when x"47B" => data <= "0111000111";
                when x"47C" => data <= "1101010101";
                when x"47D" => data <= "0000000101";
                when x"47E" => data <= "0000000101";
                when x"47F" => data <= "1100111111";
                when x"480" => data <= "1100111111";
                when x"481" => data <= "1111101011";
                when x"482" => data <= "0000000101";
                when x"483" => data <= "1011111101";
                when x"484" => data <= "0000000101";
                when x"485" => data <= "0001011010";
                when x"486" => data <= "1011111101";
                when x"487" => data <= "0000000101";
                when x"488" => data <= "1011001000";
                when x"489" => data <= "0001000000";
                when x"48A" => data <= "0100001001";
                when x"48B" => data <= "0001000000";
                when x"48C" => data <= "1011010010";
                when x"48D" => data <= "0111011101";
                when x"48E" => data <= "1011100111";
                when x"48F" => data <= "0101010110";
                when x"490" => data <= "1101111010";
                when x"491" => data <= "0110000010";
                when x"492" => data <= "0001000000";
                when x"493" => data <= "0001000000";
                when x"494" => data <= "1011010010";
                when x"495" => data <= "0001000000";
                when x"496" => data <= "0001110101";
                when x"497" => data <= "0001000000";
                when x"498" => data <= "1011010010";
                when x"499" => data <= "0001000000";
                when x"49A" => data <= "0011001011";
                when x"49B" => data <= "1110101110";
                when x"49C" => data <= "1100010000";
                when x"49D" => data <= "0110000010";
                when x"49E" => data <= "1010111000";
                when x"49F" => data <= "0110000010";
                when x"4A0" => data <= "0001000000";
                when x"4A1" => data <= "0001000000";
                when x"4A2" => data <= "0010100001";
                when x"4A3" => data <= "1000110011";
                when x"4A4" => data <= "0001000000";
                when x"4A5" => data <= "1000110011";
                when x"4A6" => data <= "0001000000";
                when x"4A7" => data <= "0001000000";
                when x"4A8" => data <= "0001000000";
                when x"4A9" => data <= "0111101000";
                when x"4AA" => data <= "0001000000";
                when x"4AB" => data <= "1100010000";
                when x"4AC" => data <= "0001000000";
                when x"4AD" => data <= "0001000000";
                when x"4AE" => data <= "0100001001";
                when x"4AF" => data <= "0110000010";
                when x"4B0" => data <= "1111000100";
                when x"4B1" => data <= "0001000000";
                when x"4B2" => data <= "1011100111";
                when x"4B3" => data <= "0001000000";
                when x"4B4" => data <= "1011100111";
                when x"4B5" => data <= "0001000000";
                when x"4B6" => data <= "0001000000";
                when x"4B7" => data <= "0001000000";
                when x"4B8" => data <= "0001000000";
                when x"4B9" => data <= "0001000000";
                when x"4BA" => data <= "0001000000";
                when x"4BB" => data <= "0001000000";
                when x"4BC" => data <= "1010111000";
                when x"4BD" => data <= "0001000000";
                when x"4BE" => data <= "1011100111";
                when x"4BF" => data <= "1100100101";
                when x"4C0" => data <= "0001000000";
                when x"4C1" => data <= "0001000000";
                when x"4C2" => data <= "0001000000";
                when x"4C3" => data <= "1011100111";
                when x"4C4" => data <= "0000101010";
                when x"4C5" => data <= "0111101000";
                when x"4C6" => data <= "0001000000";
                when x"4C7" => data <= "0110110111";
                when x"4C8" => data <= "1011100111";
                when x"4C9" => data <= "0001000000";
                when x"4CA" => data <= "0001000000";
                when x"4CB" => data <= "0111101000";
                when x"4CC" => data <= "1001011001";
                when x"4CD" => data <= "1111000100";
                when x"4CE" => data <= "0111111111";
                when x"4CF" => data <= "0000001000";
                when x"4D0" => data <= "0111111111";
                when x"4D1" => data <= "0000001000";
                when x"4D2" => data <= "1000100100";
                when x"4D3" => data <= "1010101111";
                when x"4D4" => data <= "0111111111";
                when x"4D5" => data <= "1011000101";
                when x"4D6" => data <= "0000001000";
                when x"4D7" => data <= "0111111111";
                when x"4D8" => data <= "0111111111";
                when x"4D9" => data <= "0000001000";
                when x"4DA" => data <= "0111111111";
                when x"4DB" => data <= "0000001000";
                when x"4DC" => data <= "0000001000";
                when x"4DD" => data <= "0000001000";
                when x"4DE" => data <= "1001111011";
                when x"4DF" => data <= "0111111111";
                when x"4E0" => data <= "0111111111";
                when x"4E1" => data <= "1010101111";
                when x"4E2" => data <= "0111111111";
                when x"4E3" => data <= "0111001010";
                when x"4E4" => data <= "0111111111";
                when x"4E5" => data <= "0111111111";
                when x"4E6" => data <= "0000111101";
                when x"4E7" => data <= "0111111111";
                when x"4E8" => data <= "0000001000";
                when x"4E9" => data <= "0111111111";
                when x"4EA" => data <= "0111111111";
                when x"4EB" => data <= "0111111111";
                when x"4EC" => data <= "0111111111";
                when x"4ED" => data <= "0000001000";
                when x"4EE" => data <= "0111111111";
                when x"4EF" => data <= "0111111111";
                when x"4F0" => data <= "0111111111";
                when x"4F1" => data <= "0111111111";
                when x"4F2" => data <= "0111111111";
                when x"4F3" => data <= "0111111111";
                when x"4F4" => data <= "0111111111";
                when x"4F5" => data <= "1110111001";
                when x"4F6" => data <= "1010101111";
                when x"4F7" => data <= "0111111111";
                when x"4F8" => data <= "0111111111";
                when x"4F9" => data <= "0111111111";
                when x"4FA" => data <= "0000001000";
                when x"4FB" => data <= "0111111111";
                when x"4FC" => data <= "1000010001";
                when x"4FD" => data <= "0111111111";
                when x"4FE" => data <= "0000001000";
                when x"4FF" => data <= "0111111111";
                when x"500" => data <= "1001111011";
                when x"501" => data <= "0000001000";
                when x"502" => data <= "0000001000";
                when x"503" => data <= "1001111011";
                when x"504" => data <= "0000001000";
                when x"505" => data <= "0111111111";
                when x"506" => data <= "0111111111";
                when x"507" => data <= "1010101111";
                when x"508" => data <= "0000001000";
                when x"509" => data <= "0111111111";
                when x"50A" => data <= "0111111111";
                when x"50B" => data <= "0111111111";
                when x"50C" => data <= "1010101111";
                when x"50D" => data <= "0000001000";
                when x"50E" => data <= "0111111111";
                when x"50F" => data <= "0111111111";
                when x"510" => data <= "0111111111";
                when x"511" => data <= "0111111111";
                when x"512" => data <= "0111111111";
                when x"513" => data <= "0111111111";
                when x"514" => data <= "0111111111";
                when x"515" => data <= "1001111011";
                when x"516" => data <= "0000001000";
                when x"517" => data <= "1010101111";
                when x"518" => data <= "0111111111";
                when x"519" => data <= "0111111111";
                when x"51A" => data <= "0111111111";
                when x"51B" => data <= "0111111111";
                when x"51C" => data <= "0111111111";
                when x"51D" => data <= "0111111111";
                when x"51E" => data <= "0001010111";
                when x"51F" => data <= "0110100000";
                when x"520" => data <= "0111111111";
                when x"521" => data <= "0111111111";
                when x"522" => data <= "0111111111";
                when x"523" => data <= "0000001000";
                when x"524" => data <= "0111111111";
                when x"525" => data <= "0111111111";
                when x"526" => data <= "0111111111";
                when x"527" => data <= "1010101111";
                when x"528" => data <= "0111111111";
                when x"529" => data <= "0000001000";
                when x"52A" => data <= "0111111111";
                when x"52B" => data <= "0111111111";
                when x"52C" => data <= "0111111111";
                when x"52D" => data <= "0011101001";
                when x"52E" => data <= "0111111111";
                when x"52F" => data <= "0001010111";
                when x"530" => data <= "1001111011";
                when x"531" => data <= "0111001010";
                when x"532" => data <= "0000001000";
                when x"533" => data <= "0111111111";
                when x"534" => data <= "0111111111";
                when x"535" => data <= "0111111111";
                when x"536" => data <= "0000001000";
                when x"537" => data <= "0111111111";
                when x"538" => data <= "0111111111";
                when x"539" => data <= "0111111111";
                when x"53A" => data <= "0111111111";
                when x"53B" => data <= "0111111111";
                when x"53C" => data <= "0111111111";
                when x"53D" => data <= "0111111111";
                when x"53E" => data <= "0111111111";
                when x"53F" => data <= "0111111111";
                when x"540" => data <= "0000001000";
                when x"541" => data <= "0111111111";
                when x"542" => data <= "0111111111";
                when x"543" => data <= "0111111111";
                when x"544" => data <= "0111111111";
                when x"545" => data <= "0111111111";
                when x"546" => data <= "1010011010";
                when x"547" => data <= "0111111111";
                when x"548" => data <= "0111111111";
                when x"549" => data <= "0111111111";
                when x"54A" => data <= "0111111111";
                when x"54B" => data <= "0111111111";
                when x"54C" => data <= "0111111111";
                when x"54D" => data <= "0111111111";
                when x"54E" => data <= "0111111111";
                when x"54F" => data <= "0110100000";
                when x"550" => data <= "1000100100";
                when x"551" => data <= "1110111001";
                when x"552" => data <= "0111111111";
                when x"553" => data <= "0000001000";
                when x"554" => data <= "1010101111";
                when x"555" => data <= "0000001000";
                when x"556" => data <= "0111111111";
                when x"557" => data <= "0111111111";
                when x"558" => data <= "0111111111";
                when x"559" => data <= "0111111111";
                when x"55A" => data <= "0111111111";
                when x"55B" => data <= "0111111111";
                when x"55C" => data <= "0111111111";
                when x"55D" => data <= "0111111111";
                when x"55E" => data <= "0111111111";
                when x"55F" => data <= "0111111111";
                when x"560" => data <= "0111111111";
                when x"561" => data <= "0000001000";
                when x"562" => data <= "0000001000";
                when x"563" => data <= "0000001000";
                when x"564" => data <= "0111111111";
                when x"565" => data <= "0111111111";
                when x"566" => data <= "0111111111";
                when x"567" => data <= "0000001000";
                when x"568" => data <= "0000001000";
                when x"569" => data <= "0000001000";
                when x"56A" => data <= "0111111111";
                when x"56B" => data <= "0111111111";
                when x"56C" => data <= "0000001000";
                when x"56D" => data <= "0111111111";
                when x"56E" => data <= "0111111111";
                when x"56F" => data <= "0000001000";
                when x"570" => data <= "0111111111";
                when x"571" => data <= "0111111111";
                when x"572" => data <= "0000001000";
                when x"573" => data <= "0111111111";
                when x"574" => data <= "0000001000";
                when x"575" => data <= "0111111111";
                when x"576" => data <= "0111111111";
                when x"577" => data <= "0111111111";
                when x"578" => data <= "1001111011";
                when x"579" => data <= "0001010111";
                when x"57A" => data <= "0111111111";
                when x"57B" => data <= "0111111111";
                when x"57C" => data <= "0111111111";
                when x"57D" => data <= "0111111111";
                when x"57E" => data <= "0111111111";
                when x"57F" => data <= "1010011010";
                when x"580" => data <= "0111111111";
                when x"581" => data <= "0111111111";
                when x"582" => data <= "0000001000";
                when x"583" => data <= "0111111111";
                when x"584" => data <= "0000001000";
                when x"585" => data <= "0000001000";
                when x"586" => data <= "0111111111";
                when x"587" => data <= "0111111111";
                when x"588" => data <= "0111111111";
                when x"589" => data <= "0111111111";
                when x"58A" => data <= "0111111111";
                when x"58B" => data <= "0000010010";
                when x"58C" => data <= "0000010010";
                when x"58D" => data <= "1010000000";
                when x"58E" => data <= "1010000000";
                when x"58F" => data <= "0000100111";
                when x"590" => data <= "0000100111";
                when x"591" => data <= "1101110111";
                when x"592" => data <= "0110111010";
                when x"593" => data <= "1101110111";
                when x"594" => data <= "1101110111";
                when x"595" => data <= "1101110111";
                when x"596" => data <= "0111100101";
                when x"597" => data <= "0100000100";
                when x"598" => data <= "1010000000";
                when x"599" => data <= "1101110111";
                when x"59A" => data <= "1100101000";
                when x"59B" => data <= "1101110111";
                when x"59C" => data <= "1010000000";
                when x"59D" => data <= "0111100101";
                when x"59E" => data <= "0100000100";
                when x"59F" => data <= "0011110011";
                when x"5A0" => data <= "1111111100";
                when x"5A1" => data <= "0111100101";
                when x"5A2" => data <= "0100000100";
                when x"5A3" => data <= "0110111010";
                when x"5A4" => data <= "1011011111";
                when x"5A5" => data <= "0100000100";
                when x"5A6" => data <= "1101110111";
                when x"5A7" => data <= "1101110111";
                when x"5A8" => data <= "0100000100";
                when x"5A9" => data <= "1100011101";
                when x"5AA" => data <= "0011000110";
                when x"5AB" => data <= "1101110111";
                when x"5AC" => data <= "0010101100";
                when x"5AD" => data <= "1011011111";
                when x"5AE" => data <= "0100000100";
                when x"5AF" => data <= "1011011111";
                when x"5B0" => data <= "0100000100";
                when x"5B1" => data <= "1101110111";
                when x"5B2" => data <= "1100101000";
                when x"5B3" => data <= "0100000100";
                when x"5B4" => data <= "0111010000";
                when x"5B5" => data <= "1010000000";
                when x"5B6" => data <= "0111100101";
                when x"5B7" => data <= "1010000000";
                when x"5B8" => data <= "0100000100";
                when x"5B9" => data <= "0101011011";
                when x"5BA" => data <= "1010000000";
                when x"5BB" => data <= "0100000100";
                when x"5BC" => data <= "1100011101";
                when x"5BD" => data <= "1010000000";
                when x"5BE" => data <= "1101110111";
                when x"5BF" => data <= "1010000000";
                when x"5C0" => data <= "0100000100";
                when x"5C1" => data <= "1001010100";
                when x"5C2" => data <= "1010000000";
                when x"5C3" => data <= "1010000000";
                when x"5C4" => data <= "0010101100";
                when x"5C5" => data <= "0100000100";
                when x"5C6" => data <= "1101110111";
                when x"5C7" => data <= "1100011101";
                when x"5C8" => data <= "1101110111";
                when x"5C9" => data <= "1011011111";
                when x"5CA" => data <= "1101000010";
                when x"5CB" => data <= "0110111010";
                when x"5CC" => data <= "1101110111";
                when x"5CD" => data <= "0100000100";
                when x"5CE" => data <= "1000110101";
                when x"5CF" => data <= "1111110111";
                when x"5D0" => data <= "1000000000";
                when x"5D1" => data <= "1111110111";
                when x"5D2" => data <= "1111110111";
                when x"5D3" => data <= "1111110111";
                when x"5D4" => data <= "1000000000";
                when x"5D5" => data <= "1000000000";
                when x"5D6" => data <= "1000000000";
                when x"5D7" => data <= "1111110111";
                when x"5D8" => data <= "1000000000";
                when x"5D9" => data <= "1000000000";
                when x"5DA" => data <= "1000000000";
                when x"5DB" => data <= "1000000000";
                when x"5DC" => data <= "1000000000";
                when x"5DD" => data <= "1111110111";
                when x"5DE" => data <= "1000000000";
                when x"5DF" => data <= "1111110111";
                when x"5E0" => data <= "1010111110";
                when x"5E1" => data <= "1000000000";
                when x"5E2" => data <= "1000000000";
                when x"5E3" => data <= "0110000100";
                when x"5E4" => data <= "1000000000";
                when x"5E5" => data <= "1000000000";
                when x"5E6" => data <= "1000000000";
                when x"5E7" => data <= "1111110111";
                when x"5E8" => data <= "1000000000";
                when x"5E9" => data <= "1000110101";
                when x"5EA" => data <= "1000000000";
                when x"5EB" => data <= "1000000000";
                when x"5EC" => data <= "1000000000";
                when x"5ED" => data <= "1111110111";
                when x"5EE" => data <= "1111110111";
                when x"5EF" => data <= "1000000000";
                when x"5F0" => data <= "1111110111";
                when x"5F1" => data <= "1000000000";
                when x"5F2" => data <= "1000000000";
                when x"5F3" => data <= "1000000000";
                when x"5F4" => data <= "1111110111";
                when x"5F5" => data <= "1000000000";
                when x"5F6" => data <= "1000000000";
                when x"5F7" => data <= "1000000000";
                when x"5F8" => data <= "1000000000";
                when x"5F9" => data <= "1000110101";
                when x"5FA" => data <= "1000000000";
                when x"5FB" => data <= "1000000000";
                when x"5FC" => data <= "0111011011";
                when x"5FD" => data <= "1000000000";
                when x"5FE" => data <= "1000000000";
                when x"5FF" => data <= "0101100101";
                when x"600" => data <= "1111110111";
                when x"601" => data <= "1000000000";
                when x"602" => data <= "1000000000";
                when x"603" => data <= "1000000000";
                when x"604" => data <= "1111110111";
                when x"605" => data <= "1110101000";
                when x"606" => data <= "1000000000";
                when x"607" => data <= "1000000000";
                when x"608" => data <= "1111110111";
                when x"609" => data <= "1000000000";
                when x"60A" => data <= "1000000000";
                when x"60B" => data <= "1111110111";
                when x"60C" => data <= "1111110111";
                when x"60D" => data <= "1000000000";
                when x"60E" => data <= "1000000000";
                when x"60F" => data <= "1001011111";
                when x"610" => data <= "1111110111";
                when x"611" => data <= "1011100001";
                when x"612" => data <= "1000000000";
                when x"613" => data <= "1000000000";
                when x"614" => data <= "1111000010";
                when x"615" => data <= "0000101100";
                when x"616" => data <= "1000000000";
                when x"617" => data <= "1111110111";
                when x"618" => data <= "0101010000";
                when x"619" => data <= "1111110111";
                when x"61A" => data <= "1000000000";
                when x"61B" => data <= "1000000000";
                when x"61C" => data <= "1111110111";
                when x"61D" => data <= "1110101000";
                when x"61E" => data <= "1000000000";
                when x"61F" => data <= "1000000000";
                when x"620" => data <= "1000000000";
                when x"621" => data <= "1000000000";
                when x"622" => data <= "1000000000";
                when x"623" => data <= "1000000000";
                when x"624" => data <= "1000110101";
                when x"625" => data <= "1000000000";
                when x"626" => data <= "1000000000";
                when x"627" => data <= "1111110111";
                when x"628" => data <= "1000000000";
                when x"629" => data <= "1111110111";
                when x"62A" => data <= "1000000000";
                when x"62B" => data <= "1000000000";
                when x"62C" => data <= "1000000000";
                when x"62D" => data <= "1111110111";
                when x"62E" => data <= "1000000000";
                when x"62F" => data <= "1000000000";
                when x"630" => data <= "1000000000";
                when x"631" => data <= "1000000000";
                when x"632" => data <= "1111110111";
                when x"633" => data <= "1000000000";
                when x"634" => data <= "1000000000";
                when x"635" => data <= "1000000000";
                when x"636" => data <= "1111110111";
                when x"637" => data <= "1000000000";
                when x"638" => data <= "1111110111";
                when x"639" => data <= "1000000000";
                when x"63A" => data <= "1000000000";
                when x"63B" => data <= "0110000100";
                when x"63C" => data <= "1111110111";
                when x"63D" => data <= "1000000000";
                when x"63E" => data <= "1111110111";
                when x"63F" => data <= "1000000000";
                when x"640" => data <= "0101100101";
                when x"641" => data <= "1000000000";
                when x"642" => data <= "1000000000";
                when x"643" => data <= "1000000000";
                when x"644" => data <= "1000000000";
                when x"645" => data <= "0001110011";
                when x"646" => data <= "1000000000";
                when x"647" => data <= "1000000000";
                when x"648" => data <= "1000000000";
                when x"649" => data <= "1000000000";
                when x"64A" => data <= "1000000000";
                when x"64B" => data <= "1000000000";
                when x"64C" => data <= "1111110111";
                when x"64D" => data <= "1000000000";
                when x"64E" => data <= "0101010000";
                when x"64F" => data <= "1000000000";
                when x"650" => data <= "1000000000";
                when x"651" => data <= "1000000000";
                when x"652" => data <= "1000000000";
                when x"653" => data <= "1111110111";
                when x"654" => data <= "1000000000";
                when x"655" => data <= "1000000000";
                when x"656" => data <= "0101010000";
                when x"657" => data <= "1000000000";
                when x"658" => data <= "0101010000";
                when x"659" => data <= "1000110101";
                when x"65A" => data <= "1000000000";
                when x"65B" => data <= "1111110111";
                when x"65C" => data <= "1111110111";
                when x"65D" => data <= "1111110111";
                when x"65E" => data <= "1000000000";
                when x"65F" => data <= "0101010000";
                when x"660" => data <= "1111110111";
                when x"661" => data <= "0101010000";
                when x"662" => data <= "1000000000";
                when x"663" => data <= "1111110111";
                when x"664" => data <= "1000000000";
                when x"665" => data <= "1111110111";
                when x"666" => data <= "1111110111";
                when x"667" => data <= "1111110111";
                when x"668" => data <= "1111110111";
                when x"669" => data <= "1000000000";
                when x"66A" => data <= "1000000000";
                when x"66B" => data <= "1111110111";
                when x"66C" => data <= "1000000000";
                when x"66D" => data <= "1000000000";
                when x"66E" => data <= "1000000000";
                when x"66F" => data <= "1000000000";
                when x"670" => data <= "1000000000";
                when x"671" => data <= "1000000000";
                when x"672" => data <= "1111110111";
                when x"673" => data <= "1000000000";
                when x"674" => data <= "1000000000";
                when x"675" => data <= "0101100101";
                when x"676" => data <= "1000000000";
                when x"677" => data <= "0101100101";
                when x"678" => data <= "1111110111";
                when x"679" => data <= "1000000000";
                when x"67A" => data <= "1111110111";
                when x"67B" => data <= "1110101000";
                when x"67C" => data <= "1000000000";
                when x"67D" => data <= "1000000000";
                when x"67E" => data <= "1111110111";
                when x"67F" => data <= "1000000000";
                when x"680" => data <= "1111110111";
                when x"681" => data <= "1000000000";
                when x"682" => data <= "1000000000";
                when x"683" => data <= "1000000000";
                when x"684" => data <= "1000000000";
                when x"685" => data <= "1000000000";
                when x"686" => data <= "1111110111";
                when x"687" => data <= "1000000000";
                when x"688" => data <= "1111110111";
                when x"689" => data <= "1011010100";
                when x"68A" => data <= "1000000000";
                when x"68B" => data <= "1111110111";
                when x"68C" => data <= "1111110111";
                when x"68D" => data <= "0101010000";
                when x"68E" => data <= "1000000000";
                when x"68F" => data <= "1111110111";
                when x"690" => data <= "1000000000";
                when x"691" => data <= "1000000000";
                when x"692" => data <= "0010001000";
                when x"693" => data <= "0101111111";
                when x"694" => data <= "0101111111";
                when x"695" => data <= "1011111011";
                when x"696" => data <= "1111101101";
                when x"697" => data <= "0101111111";
                when x"698" => data <= "0100100000";
                when x"699" => data <= "1011111011";
                when x"69A" => data <= "0010001000";
                when x"69B" => data <= "0101111111";
                when x"69C" => data <= "1011111011";
                when x"69D" => data <= "0100010101";
                when x"69E" => data <= "0101111111";
                when x"69F" => data <= "0100010101";
                when x"6A0" => data <= "1111011000";
                when x"6A1" => data <= "0101001010";
                when x"6A2" => data <= "0010001000";
                when x"6A3" => data <= "1011111011";
                when x"6A4" => data <= "0010001000";
                when x"6A5" => data <= "0001101001";
                when x"6A6" => data <= "0010001000";
                when x"6A7" => data <= "1011111011";
                when x"6A8" => data <= "1111011000";
                when x"6A9" => data <= "0010001000";
                when x"6AA" => data <= "0010001000";
                when x"6AB" => data <= "0100010101";
                when x"6AC" => data <= "1111011000";
                when x"6AD" => data <= "1011111011";
                when x"6AE" => data <= "0010001000";
                when x"6AF" => data <= "1011111011";
                when x"6B0" => data <= "0010001000";
                when x"6B1" => data <= "1001110000";
                when x"6B2" => data <= "1011111011";
                when x"6B3" => data <= "1011111011";
                when x"6B4" => data <= "0100100000";
                when x"6B5" => data <= "0010001000";
                when x"6B6" => data <= "1011111011";
                when x"6B7" => data <= "0101111111";
                when x"6B8" => data <= "1111011000";
                when x"6B9" => data <= "0101111111";
                when x"6BA" => data <= "1011111011";
                when x"6BB" => data <= "0010001000";
                when x"6BC" => data <= "1011111011";
                when x"6BD" => data <= "1101010011";
                when x"6BE" => data <= "0000000011";
                when x"6BF" => data <= "1111011000";
                when x"6C0" => data <= "0010001000";
                when x"6C1" => data <= "0010001000";
                when x"6C2" => data <= "1011111011";
                when x"6C3" => data <= "1011111011";
                when x"6C4" => data <= "0010001000";
                when x"6C5" => data <= "1011111011";
                when x"6C6" => data <= "0101111111";
                when x"6C7" => data <= "0100100000";
                when x"6C8" => data <= "0101111111";
                when x"6C9" => data <= "1011111011";
                when x"6CA" => data <= "0010001000";
                when x"6CB" => data <= "1111011000";
                when x"6CC" => data <= "0101111111";
                when x"6CD" => data <= "0010001000";
                when x"6CE" => data <= "0101111111";
                when x"6CF" => data <= "1011111011";
                when x"6D0" => data <= "0100100000";
                when x"6D1" => data <= "0101111111";
                when x"6D2" => data <= "0101111111";
                when x"6D3" => data <= "1011001110";
                when x"6D4" => data <= "0101111111";
                when x"6D5" => data <= "0010001000";
                when x"6D6" => data <= "0110101011";
                when x"6D7" => data <= "1000101111";
                when x"6D8" => data <= "0101111111";
                when x"6D9" => data <= "1011111011";
                when x"6DA" => data <= "1011111011";
                when x"6DB" => data <= "0010001000";
                when x"6DC" => data <= "0101111111";
                when x"6DD" => data <= "1011111011";
                when x"6DE" => data <= "0010101010";
                when x"6DF" => data <= "0100110111";
                when x"6E0" => data <= "1001010010";
                when x"6E1" => data <= "1111111010";
                when x"6E2" => data <= "1111111010";
                when x"6E3" => data <= "0100000010";
                when x"6E4" => data <= "1010110011";
                when x"6E5" => data <= "0000100001";
                when x"6E6" => data <= "1111111010";
                when x"6E7" => data <= "0100000010";
                when x"6E8" => data <= "0011000000";
                when x"6E9" => data <= "1000111000";
                when x"6EA" => data <= "1001010010";
                when x"6EB" => data <= "0000100001";
                when x"6EC" => data <= "1001010010";
                when x"6ED" => data <= "0100000010";
                when x"6EE" => data <= "0110111100";
                when x"6EF" => data <= "1001010010";
                when x"6F0" => data <= "0000100001";
                when x"6F1" => data <= "0011000000";
                when x"6F2" => data <= "1111111010";
                when x"6F3" => data <= "1111111010";
                when x"6F4" => data <= "0010101010";
                when x"6F5" => data <= "0001001011";
                when x"6F6" => data <= "1011011001";
                when x"6F7" => data <= "0111010110";
                when x"6F8" => data <= "1001010010";
                when x"6F9" => data <= "1001010010";
                when x"6FA" => data <= "0111010110";
                when x"6FB" => data <= "0100110111";
                when x"6FC" => data <= "1000111000";
                when x"6FD" => data <= "0011000000";
                when x"6FE" => data <= "1000111000";
                when x"6FF" => data <= "1111001111";
                when x"700" => data <= "1111111010";
                when x"701" => data <= "0001001011";
                when x"702" => data <= "0100110111";
                when x"703" => data <= "0011000000";
                when x"704" => data <= "1111111010";
                when x"705" => data <= "1111111010";
                when x"706" => data <= "0101011101";
                when x"707" => data <= "1111111010";
                when x"708" => data <= "0000100001";
                when x"709" => data <= "1001010010";
                when x"70A" => data <= "1001010010";
                when x"70B" => data <= "1000001101";
                when x"70C" => data <= "0100000010";
                when x"70D" => data <= "0011000000";
                when x"70E" => data <= "0100000010";
                when x"70F" => data <= "1000111000";
                when x"710" => data <= "0111010110";
                when x"711" => data <= "0101011101";
                when x"712" => data <= "0011000000";
                when x"713" => data <= "0000100001";
                when x"714" => data <= "1111111010";
                when x"715" => data <= "0000100001";
                when x"716" => data <= "1111111010";
                when x"717" => data <= "0001111110";
                when x"718" => data <= "1111111010";
                when x"719" => data <= "1000001101";
                when x"71A" => data <= "1111111010";
                when x"71B" => data <= "0000010100";
                when x"71C" => data <= "1101110001";
                when x"71D" => data <= "1000111000";
                when x"71E" => data <= "0000100001";
                when x"71F" => data <= "1111111010";
                when x"720" => data <= "1000111000";
                when x"721" => data <= "0100000010";
                when x"722" => data <= "0100000010";
                when x"723" => data <= "1111111010";
                when x"724" => data <= "1001001000";
                when x"725" => data <= "0010000101";
                when x"726" => data <= "1110111111";
                when x"727" => data <= "1010101001";
                when x"728" => data <= "0000111011";
                when x"729" => data <= "0111001100";
                when x"72A" => data <= "0011101111";
                when x"72B" => data <= "0001100100";
                when x"72C" => data <= "0100101101";
                when x"72D" => data <= "1110111111";
                when x"72E" => data <= "0011011010";
                when x"72F" => data <= "1110111111";
                when x"730" => data <= "1110111111";
                when x"731" => data <= "1110111111";
                when x"732" => data <= "1110111111";
                when x"733" => data <= "1110111111";
                when x"734" => data <= "0100101101";
                when x"735" => data <= "1001111101";
                when x"736" => data <= "0010000101";
                when x"737" => data <= "0010000101";
                when x"738" => data <= "1101011110";
                when x"739" => data <= "1110111111";
                when x"73A" => data <= "1110111111";
                when x"73B" => data <= "1110111111";
                when x"73C" => data <= "1110111111";
                when x"73D" => data <= "1110111111";
                when x"73E" => data <= "1110111111";
                when x"73F" => data <= "1001111101";
                when x"740" => data <= "0100101101";
                when x"741" => data <= "1100110100";
                when x"742" => data <= "1110111111";
                when x"743" => data <= "1110111111";
                when x"744" => data <= "1110111111";
                when x"745" => data <= "1110111111";
                when x"746" => data <= "1001001000";
                when x"747" => data <= "1011110110";
                when x"748" => data <= "1001111101";
                when x"749" => data <= "1110111111";
                when x"74A" => data <= "0100101101";
                when x"74B" => data <= "1110111111";
                when x"74C" => data <= "1010101001";
                when x"74D" => data <= "1110111111";
                when x"74E" => data <= "1110111111";
                when x"74F" => data <= "0100101101";
                when x"750" => data <= "0011011010";
                when x"751" => data <= "1110111111";
                when x"752" => data <= "0011101111";
                when x"753" => data <= "1001001000";
                when x"754" => data <= "1011110110";
                when x"755" => data <= "1110111111";
                when x"756" => data <= "0010000000";
                when x"757" => data <= "0010000000";
                when x"758" => data <= "0101000010";
                when x"759" => data <= "1100110001";
                when x"75A" => data <= "0010000000";
                when x"75B" => data <= "1000010010";
                when x"75C" => data <= "0010000000";
                when x"75D" => data <= "1001111000";
                when x"75E" => data <= "0010000000";
                when x"75F" => data <= "1000100111";
                when x"760" => data <= "1011000110";
                when x"761" => data <= "0010000000";
                when x"762" => data <= "0101110111";
                when x"763" => data <= "0010000000";
                when x"764" => data <= "1000100111";
                when x"765" => data <= "0010000000";
                when x"766" => data <= "0010000000";
                when x"767" => data <= "0010000000";
                when x"768" => data <= "1100000100";
                when x"769" => data <= "1010101100";
                when x"76A" => data <= "0010000000";
                when x"76B" => data <= "0010000000";
                when x"76C" => data <= "0000001011";
                when x"76D" => data <= "1110111010";
                when x"76E" => data <= "0101110111";
                when x"76F" => data <= "0010000000";
                when x"770" => data <= "1111100101";
                when x"771" => data <= "1010101100";
                when x"772" => data <= "0010000000";
                when x"773" => data <= "0101110111";
                when x"774" => data <= "0101110111";
                when x"775" => data <= "0010000000";
                when x"776" => data <= "0101110111";
                when x"777" => data <= "0101000010";
                when x"778" => data <= "0101110111";
                when x"779" => data <= "1111010000";
                when x"77A" => data <= "1000010010";
                when x"77B" => data <= "1100110001";
                when x"77C" => data <= "0010000000";
                when x"77D" => data <= "0101110111";
                when x"77E" => data <= "0010000000";
                when x"77F" => data <= "0101000010";
                when x"780" => data <= "0101110111";
                when x"781" => data <= "1011110011";
                when x"782" => data <= "0010000000";
                when x"783" => data <= "1111010000";
                when x"784" => data <= "0010000000";
                when x"785" => data <= "0001010100";
                when x"786" => data <= "0010000000";
                when x"787" => data <= "0101110111";
                when x"788" => data <= "0010000000";
                when x"789" => data <= "0011101010";
                when x"78A" => data <= "1110111010";
                when x"78B" => data <= "0101000010";
                when x"78C" => data <= "0101110111";
                when x"78D" => data <= "0101000010";
                when x"78E" => data <= "0100101000";
                when x"78F" => data <= "0010000000";
                when x"790" => data <= "0010000000";
                when x"791" => data <= "0010000000";
                when x"792" => data <= "1100000100";
                when x"793" => data <= "0111111100";
                when x"794" => data <= "0010000000";
                when x"795" => data <= "0010000000";
                when x"796" => data <= "0010000000";
                when x"797" => data <= "0101110111";
                when x"798" => data <= "1000010010";
                when x"799" => data <= "0011011111";
                when x"79A" => data <= "0100101000";
                when x"79B" => data <= "0101000010";
                when x"79C" => data <= "1000010010";
                when x"79D" => data <= "0101110111";
                when x"79E" => data <= "1100000100";
                when x"79F" => data <= "0101000010";
                when x"7A0" => data <= "0010000000";
                when x"7A1" => data <= "1000100111";
                when x"7A2" => data <= "1111111111";
                when x"7A3" => data <= "1111111111";
                when x"7A4" => data <= "1111111111";
                when x"7A5" => data <= "1111111111";
                when x"7A6" => data <= "1111111111";
                when x"7A7" => data <= "1111111111";
                when x"7A8" => data <= "1111111111";
                when x"7A9" => data <= "1111111111";
                when x"7AA" => data <= "1111111111";
                when x"7AB" => data <= "1111111111";
                when x"7AC" => data <= "1111111111";
                when x"7AD" => data <= "1111111111";
                when x"7AE" => data <= "1111111111";
                when x"7AF" => data <= "1111111111";
                when x"7B0" => data <= "1111111111";
                when x"7B1" => data <= "1111111111";
                when x"7B2" => data <= "1111111111";
                when x"7B3" => data <= "1111111111";
                when x"7B4" => data <= "1111111111";
                when x"7B5" => data <= "1111111111";
                when x"7B6" => data <= "1111111111";
                when x"7B7" => data <= "1111111111";
                when x"7B8" => data <= "1111111111";
                when x"7B9" => data <= "1111111111";
                when x"7BA" => data <= "1111111111";
                when x"7BB" => data <= "1000001000";
                when x"7BC" => data <= "1111111111";
                when x"7BD" => data <= "1111111111";
                when x"7BE" => data <= "1111111111";
                when x"7BF" => data <= "1111111111";
                when x"7C0" => data <= "1111111111";
                when x"7C1" => data <= "1111111111";
                when x"7C2" => data <= "1111111111";
                when x"7C3" => data <= "1111111111";
                when x"7C4" => data <= "1111111111";
                when x"7C5" => data <= "1111111111";
                when x"7C6" => data <= "1111111111";
                when x"7C7" => data <= "1111111111";
                when x"7C8" => data <= "1111111111";
                when x"7C9" => data <= "1111111111";
                when x"7CA" => data <= "1111111111";
                when x"7CB" => data <= "1111111111";
                when x"7CC" => data <= "1111111111";
                when x"7CD" => data <= "1111111111";
                when x"7CE" => data <= "1111111111";
                when x"7CF" => data <= "1111111111";
                when x"7D0" => data <= "1111111111";
                when x"7D1" => data <= "1111111111";
                when x"7D2" => data <= "1111111111";
                when x"7D3" => data <= "1111111111";
                when x"7D4" => data <= "1111111111";
                when x"7D5" => data <= "1111111111";
                when x"7D6" => data <= "1111111111";
                when x"7D7" => data <= "1111111111";
                when x"7D8" => data <= "1111111111";
                when x"7D9" => data <= "1111111111";
                when x"7DA" => data <= "1111111111";
                when x"7DB" => data <= "1111111111";
                when x"7DC" => data <= "1111111111";
                when x"7DD" => data <= "1111111111";
                when x"7DE" => data <= "1111111111";
                when x"7DF" => data <= "1111111111";
                when x"7E0" => data <= "1111111111";
                when x"7E1" => data <= "1111111111";
                when x"7E2" => data <= "1111111111";
                when x"7E3" => data <= "1111111111";
                when x"7E4" => data <= "1111111111";
                when x"7E5" => data <= "1111111111";
                when x"7E6" => data <= "1111111111";
                when x"7E7" => data <= "1111111111";
                when x"7E8" => data <= "1111111111";
                when x"7E9" => data <= "1111111111";
                when x"7EA" => data <= "1111111111";
                when x"7EB" => data <= "1111111111";
                when x"7EC" => data <= "1111111111";
                when x"7ED" => data <= "1111111111";
                when x"7EE" => data <= "1111111111";
                when x"7EF" => data <= "1111111111";
                when x"7F0" => data <= "1111111111";
                when x"7F1" => data <= "1111111111";
                when x"7F2" => data <= "1111111111";
                when x"7F3" => data <= "1111111111";
                when x"7F4" => data <= "1111111111";
                when x"7F5" => data <= "1111111111";
                when x"7F6" => data <= "1111111111";
                when x"7F7" => data <= "1111111111";
                when x"7F8" => data <= "1111111111";
                when x"7F9" => data <= "1111111111";
                when x"7FA" => data <= "1111111111";
                when x"7FB" => data <= "1111111111";
                when x"7FC" => data <= "1111111111";
                when x"7FD" => data <= "1111111111";
                when x"7FE" => data <= "1111111111";
                when x"7FF" => data <= "1111111111";
                when x"800" => data <= "1111111111";
                when x"801" => data <= "1111111111";
                when x"802" => data <= "1111111111";
                when x"803" => data <= "1111111111";
                when x"804" => data <= "1111111111";
                when x"805" => data <= "1111111111";
                when x"806" => data <= "1111111111";
                when x"807" => data <= "1111111111";
                when x"808" => data <= "1111111111";
                when x"809" => data <= "1111111111";
                when x"80A" => data <= "1111111111";
                when x"80B" => data <= "1111111111";
                when x"80C" => data <= "1111111111";
                when x"80D" => data <= "1111111111";
                when x"80E" => data <= "1111111111";
                when x"80F" => data <= "1111111111";
                when x"810" => data <= "1111111111";
                when x"811" => data <= "1111111111";
                when x"812" => data <= "1111111111";
                when x"813" => data <= "1111111111";
                when x"814" => data <= "1111111111";
                when x"815" => data <= "1111111111";
                when x"816" => data <= "1111111111";
                when x"817" => data <= "1111111111";
                when x"818" => data <= "1111111111";
                when x"819" => data <= "1111111111";
                when x"81A" => data <= "1111111111";
                when x"81B" => data <= "1111111111";
                when x"81C" => data <= "1111111111";
                when x"81D" => data <= "1111111111";
                when x"81E" => data <= "1111111111";
                when x"81F" => data <= "1111111111";
                when x"820" => data <= "1111111111";
                when x"821" => data <= "1111111111";
                when x"822" => data <= "1111111111";
                when x"823" => data <= "1111111111";
                when x"824" => data <= "1111111111";
                when x"825" => data <= "1111111111";
                when x"826" => data <= "1111111111";
                when x"827" => data <= "1111111111";
                when x"828" => data <= "1111111111";
                when x"829" => data <= "1111111111";
                when x"82A" => data <= "1111111111";
                when x"82B" => data <= "1111111111";
                when x"82C" => data <= "1111111111";
                when x"82D" => data <= "1111111111";
                when x"82E" => data <= "1111111111";
                when x"82F" => data <= "1111111111";
                when x"830" => data <= "1111111111";
                when x"831" => data <= "1111111111";
                when x"832" => data <= "1111111111";
                when x"833" => data <= "1111111111";
                when x"834" => data <= "1111111111";
                when x"835" => data <= "1111111111";
                when x"836" => data <= "1111111111";
                when x"837" => data <= "1111111111";
                when x"838" => data <= "1111111111";
                when x"839" => data <= "1111111111";
                when x"83A" => data <= "1111111111";
                when x"83B" => data <= "1111111111";
                when x"83C" => data <= "1111111111";
                when x"83D" => data <= "1111111111";
                when x"83E" => data <= "1111111111";
                when x"83F" => data <= "1111111111";
                when x"840" => data <= "1111111111";
                when x"841" => data <= "1111111111";
                when x"842" => data <= "1111111111";
                when x"843" => data <= "1111111111";
                when x"844" => data <= "1111111111";
                when x"845" => data <= "1111111111";
                when x"846" => data <= "1111111111";
                when x"847" => data <= "1111111111";
                when x"848" => data <= "1111111111";
                when x"849" => data <= "1111111111";
                when x"84A" => data <= "1111111111";
                when x"84B" => data <= "1111111111";
                when x"84C" => data <= "1111111111";
                when x"84D" => data <= "1111111111";
                when x"84E" => data <= "1111111111";
                when x"84F" => data <= "1111111111";
                when x"850" => data <= "1111111111";
                when x"851" => data <= "1111111111";
                when x"852" => data <= "1111111111";
                when x"853" => data <= "1111111111";
                when x"854" => data <= "1111111111";
                when x"855" => data <= "1111111111";
                when x"856" => data <= "1111111111";
                when x"857" => data <= "1111111111";
                when x"858" => data <= "1111111111";
                when x"859" => data <= "1111111111";
                when x"85A" => data <= "1111111111";
                when x"85B" => data <= "1111111111";
                when x"85C" => data <= "1111111111";
                when x"85D" => data <= "1111111111";
                when x"85E" => data <= "1111111111";
                when x"85F" => data <= "1111111111";
                when x"860" => data <= "1111111111";
                when x"861" => data <= "1111111111";
                when x"862" => data <= "1111111111";
                when x"863" => data <= "1111111111";
                when x"864" => data <= "1111111111";
                when x"865" => data <= "1111111111";
                when x"866" => data <= "1111111111";
                when x"867" => data <= "1011101001";
                when x"868" => data <= "1111111111";
                when x"869" => data <= "1111111111";
                when x"86A" => data <= "1111111111";
                when x"86B" => data <= "1111111111";
                when x"86C" => data <= "1111111111";
                when x"86D" => data <= "1111111111";
                when x"86E" => data <= "1111111111";
                when x"86F" => data <= "1111111111";
                when x"870" => data <= "1111111111";
                when x"871" => data <= "1111111111";
                when x"872" => data <= "1111111111";
                when x"873" => data <= "1111111111";
                when x"874" => data <= "1111111111";
                when x"875" => data <= "1111111111";
                when x"876" => data <= "1111111111";
                when x"877" => data <= "1111111111";
                when x"878" => data <= "1111111111";
                when x"879" => data <= "1111111111";
                when x"87A" => data <= "1111111111";
                when x"87B" => data <= "1111111111";
                when x"87C" => data <= "1111111111";
                when x"87D" => data <= "1111111111";
                when x"87E" => data <= "1111111111";
                when x"87F" => data <= "1111111111";
                when x"880" => data <= "1111111111";
                when x"881" => data <= "1111111111";
                when x"882" => data <= "1111111111";
                when x"883" => data <= "1111111111";
                when x"884" => data <= "1111111111";
                when x"885" => data <= "1111111111";
                when x"886" => data <= "1111111111";
                when x"887" => data <= "1111111111";
                when x"888" => data <= "1111111111";
                when x"889" => data <= "1111111111";
                when x"88A" => data <= "1111111111";
                when x"88B" => data <= "1111111111";
                when x"88C" => data <= "1111111111";
                when x"88D" => data <= "1111111111";
                when x"88E" => data <= "1111111111";
                when x"88F" => data <= "1111111111";
                when x"890" => data <= "1111111111";
                when x"891" => data <= "1111111111";
                when x"892" => data <= "1111111111";
                when x"893" => data <= "1111111111";
                when x"894" => data <= "1111111111";
                when x"895" => data <= "1111111111";
                when x"896" => data <= "1111111111";
                when x"897" => data <= "1111111111";
                when x"898" => data <= "1111111111";
                when x"899" => data <= "1111111111";
                when x"89A" => data <= "1111111111";
                when x"89B" => data <= "1111111111";
                when x"89C" => data <= "1111111111";
                when x"89D" => data <= "1111111111";
                when x"89E" => data <= "1111111111";
                when x"89F" => data <= "1111111111";
                when x"8A0" => data <= "1111111111";
                when x"8A1" => data <= "1111111111";
                when x"8A2" => data <= "1111111111";
                when x"8A3" => data <= "1111111111";
                when x"8A4" => data <= "1111111111";
                when x"8A5" => data <= "1111111111";
                when x"8A6" => data <= "1111111111";
                when x"8A7" => data <= "1111111111";
                when x"8A8" => data <= "1111111111";
                when x"8A9" => data <= "1111111111";
                when x"8AA" => data <= "1111111111";
                when x"8AB" => data <= "1111111111";
                when x"8AC" => data <= "1111111111";
                when x"8AD" => data <= "1111111111";
                when x"8AE" => data <= "1111111111";
                when x"8AF" => data <= "1111111111";
                when x"8B0" => data <= "1111111111";
                when x"8B1" => data <= "1111111111";
                when x"8B2" => data <= "1111111111";
                when x"8B3" => data <= "1111111111";
                when x"8B4" => data <= "1111111111";
                when x"8B5" => data <= "1111111111";
                when x"8B6" => data <= "1111111111";
                when x"8B7" => data <= "1111111111";
                when x"8B8" => data <= "1111111111";
                when x"8B9" => data <= "1111111111";
                when x"8BA" => data <= "1111111111";
                when x"8BB" => data <= "1111111111";
                when x"8BC" => data <= "1111111111";
                when x"8BD" => data <= "1111111111";
                when x"8BE" => data <= "1111111111";
                when x"8BF" => data <= "1111111111";
                when x"8C0" => data <= "1111111111";
                when x"8C1" => data <= "1111111111";
                when x"8C2" => data <= "1111111111";
                when x"8C3" => data <= "1111111111";
                when x"8C4" => data <= "1111111111";
                when x"8C5" => data <= "1111111111";
                when x"8C6" => data <= "1111111111";
                when x"8C7" => data <= "1111111111";
                when x"8C8" => data <= "1111111111";
                when x"8C9" => data <= "1111111111";
                when x"8CA" => data <= "1111111111";
                when x"8CB" => data <= "1111111111";
                when x"8CC" => data <= "1111111111";
                when x"8CD" => data <= "1111111111";
                when x"8CE" => data <= "1111111111";
                when x"8CF" => data <= "1111111111";
                when x"8D0" => data <= "1111111111";
                when x"8D1" => data <= "1000001000";
                when x"8D2" => data <= "1111111111";
                when x"8D3" => data <= "1111111111";
                when x"8D4" => data <= "1111111111";
                when x"8D5" => data <= "1111111111";
                when x"8D6" => data <= "1111111111";
                when x"8D7" => data <= "1000001000";
                when x"8D8" => data <= "1111111111";
                when x"8D9" => data <= "1111111111";
                when x"8DA" => data <= "1111111111";
                when x"8DB" => data <= "1111111111";
                when x"8DC" => data <= "1111111111";
                when x"8DD" => data <= "1111111111";
                when x"8DE" => data <= "1111001010";
                when x"8DF" => data <= "1111111111";
                when x"8E0" => data <= "1111111111";
                when x"8E1" => data <= "1000001000";
                when x"8E2" => data <= "1111111111";
                when x"8E3" => data <= "1111111111";
                when x"8E4" => data <= "1111111111";
                when x"8E5" => data <= "1111111111";
                when x"8E6" => data <= "1111111111";
                when x"8E7" => data <= "1111111111";
                when x"8E8" => data <= "1111111111";
                when x"8E9" => data <= "1111111111";
                when x"8EA" => data <= "1111111111";
                when x"8EB" => data <= "1111111111";
                when x"8EC" => data <= "1111111111";
                when x"8ED" => data <= "1111111111";
                when x"8EE" => data <= "1111111111";
                when x"8EF" => data <= "1111111111";
                when x"8F0" => data <= "1111111111";
                when x"8F1" => data <= "1111111111";
                when x"8F2" => data <= "1111111111";
                when x"8F3" => data <= "1111111111";
                when x"8F4" => data <= "1111111111";
                when x"8F5" => data <= "1111111111";
                when x"8F6" => data <= "1111111111";
                when x"8F7" => data <= "1111111111";
                when x"8F8" => data <= "1111111111";
                when x"8F9" => data <= "1111111111";
                when x"8FA" => data <= "1111111111";
                when x"8FB" => data <= "1111111111";
                when x"8FC" => data <= "1111111111";
                when x"8FD" => data <= "1111111111";
                when x"8FE" => data <= "1111111111";
                when x"8FF" => data <= "1111111111";
                when x"900" => data <= "1111111111";
                when x"901" => data <= "1111111111";
                when x"902" => data <= "1111111111";
                when x"903" => data <= "1111111111";
                when x"904" => data <= "1111111111";
                when x"905" => data <= "1111111111";
                when x"906" => data <= "1111111111";
                when x"907" => data <= "1111111111";
                when x"908" => data <= "1111111111";
                when x"909" => data <= "1111111111";
                when x"90A" => data <= "1111111111";
                when x"90B" => data <= "1111111111";
                when x"90C" => data <= "1111111111";
                when x"90D" => data <= "1111111111";
                when x"90E" => data <= "1111111111";
                when x"90F" => data <= "1111111111";
                when x"910" => data <= "1111111111";
                when x"911" => data <= "1111111111";
                when x"912" => data <= "1111111111";
                when x"913" => data <= "1111111111";
                when x"914" => data <= "1111111111";
                when x"915" => data <= "1111111111";
                when x"916" => data <= "1111111111";
                when x"917" => data <= "1111111111";
                when x"918" => data <= "1111111111";
                when x"919" => data <= "1111111111";
                when x"91A" => data <= "1111111111";
                when x"91B" => data <= "1111111111";
                when x"91C" => data <= "1111111111";
                when x"91D" => data <= "1111111111";
                when x"91E" => data <= "1111111111";
                when x"91F" => data <= "1111111111";
                when x"920" => data <= "1111111111";
                when x"921" => data <= "1111111111";
                when x"922" => data <= "1111111111";
                when x"923" => data <= "1111111111";
                when x"924" => data <= "1111111111";
                when x"925" => data <= "1111111111";
                when x"926" => data <= "1111111111";
                when x"927" => data <= "1111111111";
                when x"928" => data <= "1111111111";
                when x"929" => data <= "1111111111";
                when x"92A" => data <= "1111111111";
                when x"92B" => data <= "1111111111";
                when x"92C" => data <= "1111111111";
                when x"92D" => data <= "1111111111";
                when x"92E" => data <= "1111111111";
                when x"92F" => data <= "1111111111";
                when x"930" => data <= "1111111111";
                when x"931" => data <= "1111111111";
                when x"932" => data <= "1111111111";
                when x"933" => data <= "1111111111";
                when x"934" => data <= "1111111111";
                when x"935" => data <= "1111111111";
                when x"936" => data <= "1111111111";
                when x"937" => data <= "1111111111";
                when x"938" => data <= "1111111111";
                when x"939" => data <= "1111111111";
                when x"93A" => data <= "1111111111";
                when x"93B" => data <= "1111111111";
                when x"93C" => data <= "1111111111";
                when x"93D" => data <= "1111111111";
                when x"93E" => data <= "1111111111";
                when x"93F" => data <= "1111111111";
                when x"940" => data <= "1111111111";
                when x"941" => data <= "1111111111";
                when x"942" => data <= "1111111111";
                when x"943" => data <= "1111111111";
                when x"944" => data <= "1111111111";
                when x"945" => data <= "1111111111";
                when x"946" => data <= "1111111111";
                when x"947" => data <= "1111111111";
                when x"948" => data <= "1111111111";
                when x"949" => data <= "1111111111";
                when x"94A" => data <= "1111111111";
                when x"94B" => data <= "1111111111";
                when x"94C" => data <= "1111111111";
                when x"94D" => data <= "1111111111";
                when x"94E" => data <= "1111111111";
                when x"94F" => data <= "1111111111";
                when x"950" => data <= "1111111111";
                when x"951" => data <= "1111111111";
                when x"952" => data <= "1111111111";
                when x"953" => data <= "1111111111";
                when x"954" => data <= "1111111111";
                when x"955" => data <= "1111111111";
                when x"956" => data <= "1111111111";
                when x"957" => data <= "1111111111";
                when x"958" => data <= "1111111111";
                when x"959" => data <= "1111111111";
                when x"95A" => data <= "1111111111";
                when x"95B" => data <= "1111111111";
                when x"95C" => data <= "1111111111";
                when x"95D" => data <= "1111111111";
                when x"95E" => data <= "1111111111";
                when x"95F" => data <= "1111111111";
                when x"960" => data <= "1111111111";
                when x"961" => data <= "1111111111";
                when x"962" => data <= "1111111111";
                when x"963" => data <= "1111111111";
                when x"964" => data <= "1111111111";
                when x"965" => data <= "1111111111";
                when x"966" => data <= "1111111111";
                when x"967" => data <= "1111111111";
                when x"968" => data <= "1111111111";
                when x"969" => data <= "1111111111";
                when x"96A" => data <= "1111111111";
                when x"96B" => data <= "1111111111";
                when x"96C" => data <= "1111111111";
                when x"96D" => data <= "1111111111";
                when x"96E" => data <= "1111111111";
                when x"96F" => data <= "1111111111";
                when x"970" => data <= "1111111111";
                when x"971" => data <= "1111111111";
                when x"972" => data <= "1111111111";
                when x"973" => data <= "1111111111";
                when x"974" => data <= "0010011010";
                when x"975" => data <= "1111111111";
                when x"976" => data <= "1111111111";
                when x"977" => data <= "1111111111";
                when x"978" => data <= "1111111111";
                when x"979" => data <= "1111111111";
                when x"97A" => data <= "1111111111";
                when x"97B" => data <= "1111111111";
                when x"97C" => data <= "1111111111";
                when x"97D" => data <= "1111111111";
                when x"97E" => data <= "1111111111";
                when x"97F" => data <= "1111111111";
                when x"980" => data <= "1111111111";
                when x"981" => data <= "1111111111";
                when x"982" => data <= "1111111111";
                when x"983" => data <= "1111111111";
                when x"984" => data <= "1111111111";
                when x"985" => data <= "1111111111";
                when x"986" => data <= "1111111111";
                when x"987" => data <= "1111111111";
                when x"988" => data <= "1111111111";
                when x"989" => data <= "1111111111";
                when x"98A" => data <= "1111111111";
                when x"98B" => data <= "1111111111";
                when x"98C" => data <= "1111111111";
                when x"98D" => data <= "1111111111";
                when x"98E" => data <= "1111111111";
                when x"98F" => data <= "1111111111";
                when x"990" => data <= "1111111111";
                when x"991" => data <= "1111111111";
                when x"992" => data <= "1111111111";
                when x"993" => data <= "1111111111";
                when x"994" => data <= "1111111111";
                when x"995" => data <= "1111111111";
                when x"996" => data <= "1111111111";
                when x"997" => data <= "1111111111";
                when x"998" => data <= "1111111111";
                when x"999" => data <= "1111111111";
                when x"99A" => data <= "1111111111";
                when x"99B" => data <= "1111111111";
                when x"99C" => data <= "1111111111";
                when x"99D" => data <= "1111111111";
                when x"99E" => data <= "1111111111";
                when x"99F" => data <= "1111111111";
                when x"9A0" => data <= "1111111111";
                when x"9A1" => data <= "1111111111";
                when x"9A2" => data <= "1111111111";
                when x"9A3" => data <= "1111111111";
                when x"9A4" => data <= "1111111111";
                when x"9A5" => data <= "1111111111";
                when x"9A6" => data <= "1111111111";
                when x"9A7" => data <= "1111111111";
                when x"9A8" => data <= "1111111111";
                when x"9A9" => data <= "1111111111";
                when x"9AA" => data <= "1111111111";
                when x"9AB" => data <= "1111111111";
                when x"9AC" => data <= "1111111111";
                when x"9AD" => data <= "1111111111";
                when x"9AE" => data <= "1111111111";
                when x"9AF" => data <= "1111111111";
                when x"9B0" => data <= "1111111111";
                when x"9B1" => data <= "1111111111";
                when x"9B2" => data <= "1111111111";
                when x"9B3" => data <= "1111111111";
                when x"9B4" => data <= "1111111111";
                when x"9B5" => data <= "1111111111";
                when x"9B6" => data <= "1111111111";
                when x"9B7" => data <= "1111111111";
                when x"9B8" => data <= "1111111111";
                when x"9B9" => data <= "1111111111";
                when x"9BA" => data <= "1111111111";
                when x"9BB" => data <= "1111111111";
                when x"9BC" => data <= "1111111111";
                when x"9BD" => data <= "1111111111";
                when x"9BE" => data <= "1111111111";
                when x"9BF" => data <= "1111111111";
                when x"9C0" => data <= "1111111111";
                when x"9C1" => data <= "1111111111";
                when x"9C2" => data <= "1111111111";
                when x"9C3" => data <= "1111111111";
                when x"9C4" => data <= "1111111111";
                when x"9C5" => data <= "1111111111";
                when x"9C6" => data <= "1111111111";
                when x"9C7" => data <= "1111111111";
                when x"9C8" => data <= "1111111111";
                when x"9C9" => data <= "1111111111";
                when x"9CA" => data <= "1111111111";
                when x"9CB" => data <= "1111111111";
                when x"9CC" => data <= "1111111111";
                when x"9CD" => data <= "1111111111";
                when x"9CE" => data <= "1111111111";
                when x"9CF" => data <= "1111111111";
                when x"9D0" => data <= "1111111111";
                when x"9D1" => data <= "1111111111";
                when x"9D2" => data <= "1111111111";
                when x"9D3" => data <= "1111111111";
                when x"9D4" => data <= "1111111111";
                when x"9D5" => data <= "1111111111";
                when x"9D6" => data <= "1111111111";
                when x"9D7" => data <= "1111111111";
                when x"9D8" => data <= "1111111111";
                when x"9D9" => data <= "1111111111";
                when x"9DA" => data <= "1111111111";
                when x"9DB" => data <= "1111111111";
                when x"9DC" => data <= "1111111111";
                when x"9DD" => data <= "1111111111";
                when x"9DE" => data <= "1111111111";
                when x"9DF" => data <= "1111111111";
                when x"9E0" => data <= "1111111111";
                when x"9E1" => data <= "1111111111";
                when x"9E2" => data <= "1111111111";
                when x"9E3" => data <= "1111111111";
                when x"9E4" => data <= "1111111111";
                when x"9E5" => data <= "1111111111";
                when x"9E6" => data <= "1111111111";
                when x"9E7" => data <= "1111111111";
                when x"9E8" => data <= "1111111111";
                when x"9E9" => data <= "1111111111";
                when x"9EA" => data <= "1111111111";
                when x"9EB" => data <= "1111111111";
                when x"9EC" => data <= "1111111111";
                when x"9ED" => data <= "1111111111";
                when x"9EE" => data <= "1111111111";
                when x"9EF" => data <= "1111111111";
                when x"9F0" => data <= "1111111111";
                when x"9F1" => data <= "1111111111";
                when x"9F2" => data <= "1111111111";
                when x"9F3" => data <= "1111111111";
                when x"9F4" => data <= "1111111111";
                when x"9F5" => data <= "1111111111";
                when x"9F6" => data <= "1111111111";
                when x"9F7" => data <= "1111111111";
                when x"9F8" => data <= "1111111111";
                when x"9F9" => data <= "1111111111";
                when x"9FA" => data <= "1111111111";
                when x"9FB" => data <= "1111111111";
                when x"9FC" => data <= "1111111111";
                when x"9FD" => data <= "1111111111";
                when x"9FE" => data <= "1111111111";
                when x"9FF" => data <= "1111111111";
                when x"A00" => data <= "1111111111";
                when x"A01" => data <= "1111111111";
                when x"A02" => data <= "1111111111";
                when x"A03" => data <= "1111111111";
                when x"A04" => data <= "1111111111";
                when x"A05" => data <= "1111111111";
                when x"A06" => data <= "1111111111";
                when x"A07" => data <= "1111111111";
                when x"A08" => data <= "1111111111";
                when x"A09" => data <= "1111111111";
                when x"A0A" => data <= "1111111111";
                when x"A0B" => data <= "1111111111";
                when x"A0C" => data <= "1111111111";
                when x"A0D" => data <= "1111111111";
                when x"A0E" => data <= "1111111111";
                when x"A0F" => data <= "1111111111";
                when x"A10" => data <= "1111111111";
                when x"A11" => data <= "1111111111";
                when x"A12" => data <= "1111111111";
                when x"A13" => data <= "1111111111";
                when x"A14" => data <= "1111111111";
                when x"A15" => data <= "1111111111";
                when x"A16" => data <= "1111111111";
                when x"A17" => data <= "1111111111";
                when x"A18" => data <= "1111111111";
                when x"A19" => data <= "1111111111";
                when x"A1A" => data <= "1111111111";
                when x"A1B" => data <= "1111111111";
                when x"A1C" => data <= "1111111111";
                when x"A1D" => data <= "1111111111";
                when x"A1E" => data <= "1111111111";
                when x"A1F" => data <= "1111111111";
                when x"A20" => data <= "1111111111";
                when x"A21" => data <= "1111111111";
                when x"A22" => data <= "1111111111";
                when x"A23" => data <= "1111111111";
                when x"A24" => data <= "1111111111";
                when x"A25" => data <= "1111111111";
                when x"A26" => data <= "1111111111";
                when x"A27" => data <= "1111111111";
                when x"A28" => data <= "1111111111";
                when x"A29" => data <= "1111111111";
                when x"A2A" => data <= "1111111111";
                when x"A2B" => data <= "1111111111";
                when x"A2C" => data <= "1111111111";
                when x"A2D" => data <= "1111111111";
                when x"A2E" => data <= "1111111111";
                when x"A2F" => data <= "1111111111";
                when x"A30" => data <= "1111111111";
                when x"A31" => data <= "1111111111";
                when x"A32" => data <= "1111111111";
                when x"A33" => data <= "1111111111";
                when x"A34" => data <= "1111111111";
                when x"A35" => data <= "1111111111";
                when x"A36" => data <= "1111111111";
                when x"A37" => data <= "1111111111";
                when x"A38" => data <= "1111111111";
                when x"A39" => data <= "1111111111";
                when x"A3A" => data <= "1111111111";
                when x"A3B" => data <= "1111111111";
                when x"A3C" => data <= "1111111111";
                when x"A3D" => data <= "1111111111";
                when x"A3E" => data <= "1111111111";
                when x"A3F" => data <= "1111111111";
                when x"A40" => data <= "1111111111";
                when x"A41" => data <= "1111111111";
                when x"A42" => data <= "1111111111";
                when x"A43" => data <= "1111111111";
                when x"A44" => data <= "1111111111";
                when x"A45" => data <= "1111111111";
                when x"A46" => data <= "1111111111";
                when x"A47" => data <= "1111111111";
                when x"A48" => data <= "1111111111";
                when x"A49" => data <= "1111111111";
                when x"A4A" => data <= "1111111111";
                when x"A4B" => data <= "1111111111";
                when x"A4C" => data <= "1111111111";
                when x"A4D" => data <= "1111111111";
                when x"A4E" => data <= "1111111111";
                when x"A4F" => data <= "1111111111";
                when x"A50" => data <= "1111111111";
                when x"A51" => data <= "1111111111";
                when x"A52" => data <= "1111111111";
                when x"A53" => data <= "1111111111";
                when x"A54" => data <= "1111111111";
                when x"A55" => data <= "1111111111";
                when x"A56" => data <= "1111111111";
                when x"A57" => data <= "1111111111";
                when x"A58" => data <= "1111111111";
                when x"A59" => data <= "1111111111";
                when x"A5A" => data <= "1111111111";
                when x"A5B" => data <= "1111111111";
                when x"A5C" => data <= "1111111111";
                when x"A5D" => data <= "1111111111";
                when x"A5E" => data <= "1111111111";
                when x"A5F" => data <= "1111111111";
                when x"A60" => data <= "1111111111";
                when x"A61" => data <= "1111111111";
                when x"A62" => data <= "1111111111";
                when x"A63" => data <= "1111111111";
                when x"A64" => data <= "1111111111";
                when x"A65" => data <= "1111111111";
                when x"A66" => data <= "1111111111";
                when x"A67" => data <= "1111111111";
                when x"A68" => data <= "1111111111";
                when x"A69" => data <= "1111111111";
                when x"A6A" => data <= "1111111111";
                when x"A6B" => data <= "1111111111";
                when x"A6C" => data <= "1111111111";
                when x"A6D" => data <= "1111111111";
                when x"A6E" => data <= "1111111111";
                when x"A6F" => data <= "1111111111";
                when x"A70" => data <= "1111111111";
                when x"A71" => data <= "1111111111";
                when x"A72" => data <= "1111111111";
                when x"A73" => data <= "1111111111";
                when x"A74" => data <= "1111111111";
                when x"A75" => data <= "1111111111";
                when x"A76" => data <= "1111111111";
                when x"A77" => data <= "1111111111";
                when x"A78" => data <= "1111111111";
                when x"A79" => data <= "1111111111";
                when x"A7A" => data <= "1111111111";
                when x"A7B" => data <= "1111111111";
                when x"A7C" => data <= "1111111111";
                when x"A7D" => data <= "1111111111";
                when x"A7E" => data <= "1111111111";
                when x"A7F" => data <= "1111111111";
                when x"A80" => data <= "1111111111";
                when x"A81" => data <= "1111111111";
                when x"A82" => data <= "1111111111";
                when x"A83" => data <= "1111111111";
                when x"A84" => data <= "1111111111";
                when x"A85" => data <= "1111111111";
                when x"A86" => data <= "1111111111";
                when x"A87" => data <= "1111111111";
                when x"A88" => data <= "1111111111";
                when x"A89" => data <= "0111010011";
                when x"A8A" => data <= "1111111111";
                when x"A8B" => data <= "1111111111";
                when x"A8C" => data <= "1000001000";
                when x"A8D" => data <= "1111111111";
                when x"A8E" => data <= "1111111111";
                when x"A8F" => data <= "1111111111";
                when x"A90" => data <= "1111111111";
                when x"A91" => data <= "1111111111";
                when x"A92" => data <= "1111111111";
                when x"A93" => data <= "1111111111";
                when x"A94" => data <= "1111111111";
                when x"A95" => data <= "1111111111";
                when x"A96" => data <= "1111111111";
                when x"A97" => data <= "1111111111";
                when x"A98" => data <= "1111111111";
                when x"A99" => data <= "1111111111";
                when x"A9A" => data <= "1111111111";
                when x"A9B" => data <= "1111111111";
                when x"A9C" => data <= "1111111111";
                when x"A9D" => data <= "1111111111";
                when x"A9E" => data <= "1111111111";
                when x"A9F" => data <= "1111111111";
                when x"AA0" => data <= "1111111111";
                when x"AA1" => data <= "1111111111";
                when x"AA2" => data <= "1111111111";
                when x"AA3" => data <= "1111111111";
                when x"AA4" => data <= "1111111111";
                when x"AA5" => data <= "1111111111";
                when x"AA6" => data <= "1111111111";
                when x"AA7" => data <= "1111111111";
                when x"AA8" => data <= "1111111111";
                when x"AA9" => data <= "1111111111";
                when x"AAA" => data <= "1111111111";
                when x"AAB" => data <= "1111111111";
                when x"AAC" => data <= "1111111111";
                when x"AAD" => data <= "1111111111";
                when x"AAE" => data <= "1111111111";
                when x"AAF" => data <= "1111111111";
                when x"AB0" => data <= "1111111111";
                when x"AB1" => data <= "1111111111";
                when x"AB2" => data <= "1111111111";
                when x"AB3" => data <= "1111111111";
                when x"AB4" => data <= "1111111111";
                when x"AB5" => data <= "1111111111";
                when x"AB6" => data <= "1111111111";
                when x"AB7" => data <= "1111111111";
                when x"AB8" => data <= "1111111111";
                when x"AB9" => data <= "1111111111";
                when x"ABA" => data <= "1111111111";
                when x"ABB" => data <= "1111111111";
                when x"ABC" => data <= "1111111111";
                when x"ABD" => data <= "1111111111";
                when x"ABE" => data <= "1111111111";
                when x"ABF" => data <= "1111111111";
                when x"AC0" => data <= "1111111111";
                when x"AC1" => data <= "1111001010";
                when x"AC2" => data <= "1111111111";
                when x"AC3" => data <= "1111111111";
                when x"AC4" => data <= "1111111111";
                when x"AC5" => data <= "1111111111";
                when x"AC6" => data <= "1111111111";
                when x"AC7" => data <= "1111111111";
                when x"AC8" => data <= "1111111111";
                when x"AC9" => data <= "1111111111";
                when x"ACA" => data <= "1111111111";
                when x"ACB" => data <= "1111111111";
                when x"ACC" => data <= "1111111111";
                when x"ACD" => data <= "1111111111";
                when x"ACE" => data <= "1111111111";
                when x"ACF" => data <= "1111111111";
                when x"AD0" => data <= "1111111111";
                when x"AD1" => data <= "1111111111";
                when x"AD2" => data <= "1111111111";
                when x"AD3" => data <= "1111111111";
                when x"AD4" => data <= "1111111111";
                when x"AD5" => data <= "1111111111";
                when x"AD6" => data <= "1111111111";
                when x"AD7" => data <= "1111111111";
                when x"AD8" => data <= "1111111111";
                when x"AD9" => data <= "1111111111";
                when x"ADA" => data <= "1111111111";
                when x"ADB" => data <= "1111111111";
                when x"ADC" => data <= "1111111111";
                when x"ADD" => data <= "1111111111";
                when x"ADE" => data <= "1111111111";
                when x"ADF" => data <= "1111111111";
                when x"AE0" => data <= "1111111111";
                when x"AE1" => data <= "1111111111";
                when x"AE2" => data <= "1111111111";
                when x"AE3" => data <= "1111111111";
                when x"AE4" => data <= "1111111111";
                when x"AE5" => data <= "1111111111";
                when x"AE6" => data <= "1111111111";
                when x"AE7" => data <= "1111111111";
                when x"AE8" => data <= "1111111111";
                when x"AE9" => data <= "1111111111";
                when x"AEA" => data <= "1111111111";
                when x"AEB" => data <= "1111111111";
                when x"AEC" => data <= "1111111111";
                when x"AED" => data <= "1111111111";
                when x"AEE" => data <= "1111111111";
                when x"AEF" => data <= "1111111111";
                when x"AF0" => data <= "0010101111";
                when x"AF1" => data <= "1111111111";
                when x"AF2" => data <= "1111111111";
                when x"AF3" => data <= "1111111111";
                when x"AF4" => data <= "1111111111";
                when x"AF5" => data <= "1111111111";
                when x"AF6" => data <= "1111111111";
                when x"AF7" => data <= "1111111111";
                when x"AF8" => data <= "1111111111";
                when x"AF9" => data <= "1111111111";
                when x"AFA" => data <= "1111111111";
                when x"AFB" => data <= "1111111111";
                when x"AFC" => data <= "1111111111";
                when x"AFD" => data <= "1111111111";
                when x"AFE" => data <= "1111111111";
                when x"AFF" => data <= "1111111111";
                when x"B00" => data <= "1111111111";
                when x"B01" => data <= "1111111111";
                when x"B02" => data <= "1111111111";
                when x"B03" => data <= "1111111111";
                when x"B04" => data <= "1111111111";
                when x"B05" => data <= "1111111111";
                when x"B06" => data <= "1111111111";
                when x"B07" => data <= "1111111111";
                when x"B08" => data <= "1111111111";
                when x"B09" => data <= "1111111111";
                when x"B0A" => data <= "1111111111";
                when x"B0B" => data <= "1111111111";
                when x"B0C" => data <= "1111111111";
                when x"B0D" => data <= "1111111111";
                when x"B0E" => data <= "1111111111";
                when x"B0F" => data <= "1111111111";
                when x"B10" => data <= "1111111111";
                when x"B11" => data <= "1111111111";
                when x"B12" => data <= "1111111111";
                when x"B13" => data <= "1111111111";
                when x"B14" => data <= "1111111111";
                when x"B15" => data <= "1111111111";
                when x"B16" => data <= "1111111111";
                when x"B17" => data <= "1111111111";
                when x"B18" => data <= "1111111111";
                when x"B19" => data <= "1111111111";
                when x"B1A" => data <= "1000001000";
                when x"B1B" => data <= "1111111111";
                when x"B1C" => data <= "1111111111";
                when x"B1D" => data <= "1111111111";
                when x"B1E" => data <= "1111111111";
                when x"B1F" => data <= "1111111111";
                when x"B20" => data <= "1111111111";
                when x"B21" => data <= "1111111111";
                when x"B22" => data <= "1111111111";
                when x"B23" => data <= "1111111111";
                when x"B24" => data <= "1111111111";
                when x"B25" => data <= "1111111111";
                when x"B26" => data <= "1111111111";
                when x"B27" => data <= "1111111111";
                when x"B28" => data <= "1111111111";
                when x"B29" => data <= "1111111111";
                when x"B2A" => data <= "1111111111";
                when x"B2B" => data <= "0001111011";
                when x"B2C" => data <= "1111111111";
                when x"B2D" => data <= "1111111111";
                when x"B2E" => data <= "1111111111";
                when x"B2F" => data <= "1111111111";
                when x"B30" => data <= "1111111111";
                when x"B31" => data <= "1111111111";
                when x"B32" => data <= "1111111111";
                when x"B33" => data <= "1111111111";
                when x"B34" => data <= "1111111111";
                when x"B35" => data <= "1111111111";
                when x"B36" => data <= "1111111111";
                when x"B37" => data <= "1111111111";
                when x"B38" => data <= "1111111111";
                when x"B39" => data <= "1111111111";
                when x"B3A" => data <= "1111111111";
                when x"B3B" => data <= "1111111111";
                when x"B3C" => data <= "1111111111";
                when x"B3D" => data <= "1111111111";
                when x"B3E" => data <= "1111111111";
                when x"B3F" => data <= "1111111111";
                when x"B40" => data <= "1111111111";
                when x"B41" => data <= "1111111111";
                when x"B42" => data <= "1111111111";
                when x"B43" => data <= "1111111111";
                when x"B44" => data <= "1111111111";
                when x"B45" => data <= "1111111111";
                when x"B46" => data <= "1111111111";
                when x"B47" => data <= "1111111111";
                when x"B48" => data <= "1111111111";
                when x"B49" => data <= "1111111111";
                when x"B4A" => data <= "1111111111";
                when x"B4B" => data <= "1111111111";
                when x"B4C" => data <= "1111111111";
                when x"B4D" => data <= "1111111111";
                when x"B4E" => data <= "1111111111";
                when x"B4F" => data <= "1111111111";
                when x"B50" => data <= "1111111111";
                when x"B51" => data <= "1111111111";
                when x"B52" => data <= "1111111111";
                when x"B53" => data <= "1111111111";
                when x"B54" => data <= "1111111111";
                when x"B55" => data <= "1111111111";
                when x"B56" => data <= "1111111111";
                when x"B57" => data <= "1111111111";
                when x"B58" => data <= "1111111111";
                when x"B59" => data <= "1111111111";
                when x"B5A" => data <= "1111111111";
                when x"B5B" => data <= "1111111111";
                when x"B5C" => data <= "1111111111";
                when x"B5D" => data <= "1111111111";
                when x"B5E" => data <= "1111111111";
                when x"B5F" => data <= "1111111111";
                when x"B60" => data <= "1111111111";
                when x"B61" => data <= "1111111111";
                when x"B62" => data <= "1111111111";
                when x"B63" => data <= "1111111111";
                when x"B64" => data <= "1111111111";
                when x"B65" => data <= "1111111111";
                when x"B66" => data <= "1111111111";
                when x"B67" => data <= "1111111111";
                when x"B68" => data <= "1111111111";
                when x"B69" => data <= "1111111111";
                when x"B6A" => data <= "1111111111";
                when x"B6B" => data <= "1111111111";
                when x"B6C" => data <= "1111111111";
                when x"B6D" => data <= "1111111111";
                when x"B6E" => data <= "1111111111";
                when x"B6F" => data <= "1111111111";
                when x"B70" => data <= "1111111111";
                when x"B71" => data <= "1111111111";
                when x"B72" => data <= "1111111111";
                when x"B73" => data <= "1111111111";
                when x"B74" => data <= "1111111111";
                when x"B75" => data <= "1111111111";
                when x"B76" => data <= "1111111111";
                when x"B77" => data <= "1111111111";
                when x"B78" => data <= "1111111111";
                when x"B79" => data <= "1111111111";
                when x"B7A" => data <= "1111111111";
                when x"B7B" => data <= "1111111111";
                when x"B7C" => data <= "1111111111";
                when x"B7D" => data <= "1111111111";
                when x"B7E" => data <= "1111111111";
                when x"B7F" => data <= "1111111111";
                when x"B80" => data <= "1111111111";
                when x"B81" => data <= "1111111111";
                when x"B82" => data <= "1111111111";
                when x"B83" => data <= "1111111111";
                when x"B84" => data <= "1111111111";
                when x"B85" => data <= "1111111111";
                when x"B86" => data <= "1111111111";
                when x"B87" => data <= "1111111111";
                when x"B88" => data <= "1111111111";
                when x"B89" => data <= "1111111111";
                when x"B8A" => data <= "1111111111";
                when x"B8B" => data <= "1111111111";
                when x"B8C" => data <= "1111111111";
                when x"B8D" => data <= "1111111111";
                when x"B8E" => data <= "1111111111";
                when x"B8F" => data <= "1111111111";
                when x"B90" => data <= "1111111111";
                when x"B91" => data <= "1111111111";
                when x"B92" => data <= "1111111111";
                when x"B93" => data <= "1111111111";
                when x"B94" => data <= "1111111111";
                when x"B95" => data <= "1111111111";
                when x"B96" => data <= "1111111111";
                when x"B97" => data <= "1111111111";
                when x"B98" => data <= "1111111111";
                when x"B99" => data <= "1111111111";
                when x"B9A" => data <= "1111111111";
                when x"B9B" => data <= "1111111111";
                when x"B9C" => data <= "1111111111";
                when x"B9D" => data <= "1111111111";
                when x"B9E" => data <= "1111111111";
                when x"B9F" => data <= "1111111111";
                when x"BA0" => data <= "1111111111";
                when x"BA1" => data <= "1111111111";
                when x"BA2" => data <= "1111111111";
                when x"BA3" => data <= "1111111111";
                when x"BA4" => data <= "1111111111";
                when x"BA5" => data <= "1111111111";
                when x"BA6" => data <= "1111111111";
                when x"BA7" => data <= "1111111111";
                when x"BA8" => data <= "1111111111";
                when x"BA9" => data <= "1111111111";
                when x"BAA" => data <= "1111111111";
                when x"BAB" => data <= "1111111111";
                when x"BAC" => data <= "1111111111";
                when x"BAD" => data <= "1111111111";
                when x"BAE" => data <= "1111111111";
                when x"BAF" => data <= "1111111111";
                when x"BB0" => data <= "1111111111";
                when x"BB1" => data <= "1111111111";
                when x"BB2" => data <= "1111111111";
                when x"BB3" => data <= "1111111111";
                when x"BB4" => data <= "1111111111";
                when x"BB5" => data <= "1111111111";
                when x"BB6" => data <= "1111111111";
                when x"BB7" => data <= "1111111111";
                when x"BB8" => data <= "1111111111";
                when x"BB9" => data <= "1111111111";
                when x"BBA" => data <= "1111111111";
                when x"BBB" => data <= "1111111111";
                when x"BBC" => data <= "1111111111";
                when x"BBD" => data <= "1111111111";
                when x"BBE" => data <= "1111111111";
                when x"BBF" => data <= "1111111111";
                when x"BC0" => data <= "1111111111";
                when x"BC1" => data <= "1111111111";
                when x"BC2" => data <= "1111111111";
                when x"BC3" => data <= "1111111111";
                when x"BC4" => data <= "1111111111";
                when x"BC5" => data <= "1111111111";
                when x"BC6" => data <= "1111111111";
                when x"BC7" => data <= "1111111111";
                when x"BC8" => data <= "1111111111";
                when x"BC9" => data <= "1111111111";
                when x"BCA" => data <= "1111111111";
                when x"BCB" => data <= "1111111111";
                when x"BCC" => data <= "1111111111";
                when x"BCD" => data <= "1111111111";
                when x"BCE" => data <= "1111111111";
                when x"BCF" => data <= "1111111111";
                when x"BD0" => data <= "1111111111";
                when x"BD1" => data <= "1111111111";
                when x"BD2" => data <= "1111111111";
                when x"BD3" => data <= "1111111111";
                when x"BD4" => data <= "1111111111";
                when x"BD5" => data <= "1111111111";
                when x"BD6" => data <= "1111111111";
                when x"BD7" => data <= "1111111111";
                when x"BD8" => data <= "1111111111";
                when x"BD9" => data <= "1111111111";
                when x"BDA" => data <= "1111111111";
                when x"BDB" => data <= "1111111111";
                when x"BDC" => data <= "1111111111";
                when x"BDD" => data <= "1111111111";
                when x"BDE" => data <= "1111111111";
                when x"BDF" => data <= "1111111111";
                when x"BE0" => data <= "1111111111";
                when x"BE1" => data <= "1111111111";
                when x"BE2" => data <= "1111111111";
                when x"BE3" => data <= "1111111111";
                when x"BE4" => data <= "1111111111";
                when x"BE5" => data <= "1111111111";
                when x"BE6" => data <= "1111111111";
                when x"BE7" => data <= "1111111111";
                when x"BE8" => data <= "1111111111";
                when x"BE9" => data <= "1111111111";
                when x"BEA" => data <= "1111111111";
                when x"BEB" => data <= "1111111111";
                when x"BEC" => data <= "1001010111";
                when x"BED" => data <= "1111111111";
                when x"BEE" => data <= "1111111111";
                when x"BEF" => data <= "1111111111";
                when x"BF0" => data <= "1111111111";
                when x"BF1" => data <= "1111111111";
                when x"BF2" => data <= "1111111111";
                when x"BF3" => data <= "1111111111";
                when x"BF4" => data <= "1111111111";
                when x"BF5" => data <= "1111111111";
                when x"BF6" => data <= "1111111111";
                when x"BF7" => data <= "1111111111";
                when x"BF8" => data <= "1111111111";
                when x"BF9" => data <= "1111111111";
                when x"BFA" => data <= "1111111111";
                when x"BFB" => data <= "1111111111";
                when x"BFC" => data <= "1111111111";
                when x"BFD" => data <= "1111111111";
                when x"BFE" => data <= "1111111111";
                when x"BFF" => data <= "1111111111";
                when x"C00" => data <= "1111111111";
                when x"C01" => data <= "1111111111";
                when x"C02" => data <= "1111111111";
                when x"C03" => data <= "1111111111";
                when x"C04" => data <= "1111111111";
                when x"C05" => data <= "1111111111";
                when x"C06" => data <= "1111111111";
                when x"C07" => data <= "1111111111";
                when x"C08" => data <= "1111111111";
                when x"C09" => data <= "1111111111";
                when x"C0A" => data <= "1111111111";
                when x"C0B" => data <= "1111111111";
                when x"C0C" => data <= "1111111111";
                when x"C0D" => data <= "1111111111";
                when x"C0E" => data <= "1111111111";
                when x"C0F" => data <= "1111111111";
                when x"C10" => data <= "1111111111";
                when x"C11" => data <= "1111111111";
                when x"C12" => data <= "1111111111";
                when x"C13" => data <= "1111111111";
                when x"C14" => data <= "1111111111";
                when x"C15" => data <= "1111111111";
                when x"C16" => data <= "1111111111";
                when x"C17" => data <= "1111111111";
                when x"C18" => data <= "1111111111";
                when x"C19" => data <= "1111111111";
                when x"C1A" => data <= "1111111111";
                when x"C1B" => data <= "1111111111";
                when x"C1C" => data <= "1111111111";
                when x"C1D" => data <= "1111111111";
                when x"C1E" => data <= "1111111111";
                when x"C1F" => data <= "1111111111";
                when x"C20" => data <= "1111111111";
                when x"C21" => data <= "1111111111";
                when x"C22" => data <= "1111111111";
                when x"C23" => data <= "1111111111";
                when x"C24" => data <= "1111111111";
                when x"C25" => data <= "1111111111";
                when x"C26" => data <= "1111111111";
                when x"C27" => data <= "1111111111";
                when x"C28" => data <= "1111111111";
                when x"C29" => data <= "1111111111";
                when x"C2A" => data <= "0100000111";
                when x"C2B" => data <= "1111111111";
                when x"C2C" => data <= "1111111111";
                when x"C2D" => data <= "1111111111";
                when x"C2E" => data <= "1111111111";
                when x"C2F" => data <= "1111111111";
                when x"C30" => data <= "1111111111";
                when x"C31" => data <= "1111111111";
                when x"C32" => data <= "1111111111";
                when x"C33" => data <= "1111111111";
                when x"C34" => data <= "1111111111";
                when x"C35" => data <= "1111111111";
                when x"C36" => data <= "1111111111";
                when x"C37" => data <= "1111111111";
                when x"C38" => data <= "1111111111";
                when x"C39" => data <= "1111111111";
                when x"C3A" => data <= "1111111111";
                when x"C3B" => data <= "1111111111";
                when x"C3C" => data <= "1111111111";
                when x"C3D" => data <= "1111111111";
                when x"C3E" => data <= "1111111111";
                when x"C3F" => data <= "1111111111";
                when x"C40" => data <= "1111111111";
                when x"C41" => data <= "1111111111";
                when x"C42" => data <= "1111111111";
                when x"C43" => data <= "1111111111";
                when x"C44" => data <= "1111111111";
                when x"C45" => data <= "1111111111";
                when x"C46" => data <= "1111111111";
                when x"C47" => data <= "1111111111";
                when x"C48" => data <= "1111111111";
                when x"C49" => data <= "1111111111";
                when x"C4A" => data <= "1111111111";
                when x"C4B" => data <= "1111111111";
                when x"C4C" => data <= "1111111111";
                when x"C4D" => data <= "1111111111";
                when x"C4E" => data <= "1111111111";
                when x"C4F" => data <= "1111111111";
                when x"C50" => data <= "1111111111";
                when x"C51" => data <= "1111111111";
                when x"C52" => data <= "1111111111";
                when x"C53" => data <= "1111111111";
                when x"C54" => data <= "1111111111";
                when x"C55" => data <= "1111111111";
                when x"C56" => data <= "1111111111";
                when x"C57" => data <= "1111111111";
                when x"C58" => data <= "1111111111";
                when x"C59" => data <= "1111111111";
                when x"C5A" => data <= "1111111111";
                when x"C5B" => data <= "1111111111";
                when x"C5C" => data <= "1111111111";
                when x"C5D" => data <= "1111111111";
                when x"C5E" => data <= "1111111111";
                when x"C5F" => data <= "1111111111";
                when x"C60" => data <= "1111111111";
                when x"C61" => data <= "1111111111";
                when x"C62" => data <= "1111111111";
                when x"C63" => data <= "1111111111";
                when x"C64" => data <= "1111111111";
                when x"C65" => data <= "1111111111";
                when x"C66" => data <= "1111111111";
                when x"C67" => data <= "1111111111";
                when x"C68" => data <= "1111111111";
                when x"C69" => data <= "1111111111";
                when x"C6A" => data <= "1111111111";
                when x"C6B" => data <= "1111111111";
                when x"C6C" => data <= "1111111111";
                when x"C6D" => data <= "1111111111";
                when x"C6E" => data <= "1111111111";
                when x"C6F" => data <= "1111111111";
                when x"C70" => data <= "1111111111";
                when x"C71" => data <= "1111111111";
                when x"C72" => data <= "1111111111";
                when x"C73" => data <= "1111111111";
                when x"C74" => data <= "1111111111";
                when x"C75" => data <= "1111111111";
                when x"C76" => data <= "1111111111";
                when x"C77" => data <= "1111111111";
                when x"C78" => data <= "1111111111";
                when x"C79" => data <= "1111111111";
                when x"C7A" => data <= "1111111111";
                when x"C7B" => data <= "1111111111";
                when x"C7C" => data <= "1111111111";
                when x"C7D" => data <= "1111111111";
                when x"C7E" => data <= "1111111111";
                when x"C7F" => data <= "1111111111";
                when x"C80" => data <= "1111111111";
                when x"C81" => data <= "1111111111";
                when x"C82" => data <= "1111111111";
                when x"C83" => data <= "1111111111";
                when x"C84" => data <= "1111111111";
                when x"C85" => data <= "1111111111";
                when x"C86" => data <= "1111111111";
                when x"C87" => data <= "1111111111";
                when x"C88" => data <= "1111111111";
                when x"C89" => data <= "0001111011";
                when x"C8A" => data <= "1111111111";
                when x"C8B" => data <= "1111111111";
                when x"C8C" => data <= "1111111111";
                when x"C8D" => data <= "1111111111";
                when x"C8E" => data <= "1111111111";
                when x"C8F" => data <= "1111111111";
                when x"C90" => data <= "1111111111";
                when x"C91" => data <= "1111111111";
                when x"C92" => data <= "1111111111";
                when x"C93" => data <= "1111111111";
                when x"C94" => data <= "1111111111";
                when x"C95" => data <= "1111111111";
                when x"C96" => data <= "1111111111";
                when x"C97" => data <= "1111111111";
                when x"C98" => data <= "1111111111";
                when x"C99" => data <= "1111111111";
                when x"C9A" => data <= "1111111111";
                when x"C9B" => data <= "1111111111";
                when x"C9C" => data <= "1111111111";
                when x"C9D" => data <= "1111111111";
                when x"C9E" => data <= "1111111111";
                when x"C9F" => data <= "1111111111";
                when x"CA0" => data <= "1111111111";
                when x"CA1" => data <= "1000001000";
                when x"CA2" => data <= "1111111111";
                when x"CA3" => data <= "1111111111";
                when x"CA4" => data <= "1111111111";
                when x"CA5" => data <= "1111111111";
                when x"CA6" => data <= "1111111111";
                when x"CA7" => data <= "1111111111";
                when x"CA8" => data <= "1111111111";
                when x"CA9" => data <= "1111111111";
                when x"CAA" => data <= "1111111111";
                when x"CAB" => data <= "1111111111";
                when x"CAC" => data <= "1111111111";
                when x"CAD" => data <= "1111111111";
                when x"CAE" => data <= "1111111111";
                when x"CAF" => data <= "1111111111";
                when x"CB0" => data <= "1111111111";
                when x"CB1" => data <= "1111111111";
                when x"CB2" => data <= "1111111111";
                when x"CB3" => data <= "1111111111";
                when x"CB4" => data <= "1111111111";
                when x"CB5" => data <= "1111111111";
                when x"CB6" => data <= "1111111111";
                when x"CB7" => data <= "1111111111";
                when x"CB8" => data <= "1111111111";
                when x"CB9" => data <= "1111111111";
                when x"CBA" => data <= "1111111111";
                when x"CBB" => data <= "1111111111";
                when x"CBC" => data <= "1111111111";
                when x"CBD" => data <= "1111111111";
                when x"CBE" => data <= "1111111111";
                when x"CBF" => data <= "1111111111";
                when x"CC0" => data <= "1111111111";
                when x"CC1" => data <= "1111111111";
                when x"CC2" => data <= "1111111111";
                when x"CC3" => data <= "1111111111";
                when x"CC4" => data <= "1111111111";
                when x"CC5" => data <= "1111111111";
                when x"CC6" => data <= "1111111111";
                when x"CC7" => data <= "1111111111";
                when x"CC8" => data <= "1111111111";
                when x"CC9" => data <= "1111111111";
                when x"CCA" => data <= "1111111111";
                when x"CCB" => data <= "1111111111";
                when x"CCC" => data <= "1111111111";
                when x"CCD" => data <= "1111111111";
                when x"CCE" => data <= "1111111111";
                when x"CCF" => data <= "1111111111";
                when x"CD0" => data <= "1111111111";
                when x"CD1" => data <= "1111111111";
                when x"CD2" => data <= "1111111111";
                when x"CD3" => data <= "1111111111";
                when x"CD4" => data <= "1111111111";
                when x"CD5" => data <= "1111111111";
                when x"CD6" => data <= "1111111111";
                when x"CD7" => data <= "1111111111";
                when x"CD8" => data <= "1111111111";
                when x"CD9" => data <= "1111111111";
                when x"CDA" => data <= "1111111111";
                when x"CDB" => data <= "1111111111";
                when x"CDC" => data <= "1111111111";
                when x"CDD" => data <= "1111111111";
                when x"CDE" => data <= "1111111111";
                when x"CDF" => data <= "1111111111";
                when x"CE0" => data <= "1111111111";
                when x"CE1" => data <= "1111111111";
                when x"CE2" => data <= "1111111111";
                when x"CE3" => data <= "1111111111";
                when x"CE4" => data <= "1111111111";
                when x"CE5" => data <= "1111111111";
                when x"CE6" => data <= "1111111111";
                when x"CE7" => data <= "1111111111";
                when x"CE8" => data <= "1111111111";
                when x"CE9" => data <= "1111111111";
                when x"CEA" => data <= "1111111111";
                when x"CEB" => data <= "1111111111";
                when x"CEC" => data <= "1111111111";
                when x"CED" => data <= "1111111111";
                when x"CEE" => data <= "1111111111";
                when x"CEF" => data <= "1111111111";
                when x"CF0" => data <= "1111111111";
                when x"CF1" => data <= "1111111111";
                when x"CF2" => data <= "1111111111";
                when x"CF3" => data <= "1111111111";
                when x"CF4" => data <= "1111111111";
                when x"CF5" => data <= "1111111111";
                when x"CF6" => data <= "1111111111";
                when x"CF7" => data <= "1111111111";
                when x"CF8" => data <= "1111111111";
                when x"CF9" => data <= "1111111111";
                when x"CFA" => data <= "1111111111";
                when x"CFB" => data <= "1111111111";
                when x"CFC" => data <= "1111111111";
                when x"CFD" => data <= "1111111111";
                when x"CFE" => data <= "1111111111";
                when x"CFF" => data <= "1111111111";
                when x"D00" => data <= "1111111111";
                when x"D01" => data <= "1111111111";
                when x"D02" => data <= "1111111111";
                when x"D03" => data <= "1111111111";
                when x"D04" => data <= "1111111111";
                when x"D05" => data <= "1111111111";
                when x"D06" => data <= "1111111111";
                when x"D07" => data <= "1111111111";
                when x"D08" => data <= "1111111111";
                when x"D09" => data <= "1111111111";
                when x"D0A" => data <= "1111111111";
                when x"D0B" => data <= "1111111111";
                when x"D0C" => data <= "1111111111";
                when x"D0D" => data <= "1111111111";
                when x"D0E" => data <= "1111111111";
                when x"D0F" => data <= "1111111111";
                when x"D10" => data <= "1111111111";
                when x"D11" => data <= "1111111111";
                when x"D12" => data <= "1111111111";
                when x"D13" => data <= "1111111111";
                when x"D14" => data <= "1111111111";
                when x"D15" => data <= "1111111111";
                when x"D16" => data <= "1111111111";
                when x"D17" => data <= "1111111111";
                when x"D18" => data <= "1111111111";
                when x"D19" => data <= "1111111111";
                when x"D1A" => data <= "1111111111";
                when x"D1B" => data <= "1111111111";
                when x"D1C" => data <= "1111111111";
                when x"D1D" => data <= "1111111111";
                when x"D1E" => data <= "1111111111";
                when x"D1F" => data <= "1111111111";
                when x"D20" => data <= "1111111111";
                when x"D21" => data <= "1111111111";
                when x"D22" => data <= "1111111111";
                when x"D23" => data <= "1111111111";
                when x"D24" => data <= "1111111111";
                when x"D25" => data <= "1111111111";
                when x"D26" => data <= "1111111111";
                when x"D27" => data <= "1111111111";
                when x"D28" => data <= "1111111111";
                when x"D29" => data <= "1111111111";
                when x"D2A" => data <= "1111111111";
                when x"D2B" => data <= "1111111111";
                when x"D2C" => data <= "1111111111";
                when x"D2D" => data <= "1111111111";
                when x"D2E" => data <= "1111111111";
                when x"D2F" => data <= "1111111111";
                when x"D30" => data <= "1111111111";
                when x"D31" => data <= "1111111111";
                when x"D32" => data <= "0101011000";
                when x"D33" => data <= "1111111111";
                when x"D34" => data <= "1111111111";
                when x"D35" => data <= "1111111111";
                when x"D36" => data <= "1111111111";
                when x"D37" => data <= "1111111111";
                when x"D38" => data <= "1111111111";
                when x"D39" => data <= "1111111111";
                when x"D3A" => data <= "1111111111";
                when x"D3B" => data <= "1111111111";
                when x"D3C" => data <= "1111111111";
                when x"D3D" => data <= "1111111111";
                when x"D3E" => data <= "1111111111";
                when x"D3F" => data <= "1111111111";
                when x"D40" => data <= "1111111111";
                when x"D41" => data <= "1111111111";
                when x"D42" => data <= "1111111111";
                when x"D43" => data <= "1111111111";
                when x"D44" => data <= "1111111111";
                when x"D45" => data <= "1111111111";
                when x"D46" => data <= "1111111111";
                when x"D47" => data <= "1111111111";
                when x"D48" => data <= "1111111111";
                when x"D49" => data <= "1111111111";
                when x"D4A" => data <= "1111111111";
                when x"D4B" => data <= "1111111111";
                when x"D4C" => data <= "1111111111";
                when x"D4D" => data <= "1111111111";
                when x"D4E" => data <= "1111111111";
                when x"D4F" => data <= "1111111111";
                when x"D50" => data <= "1111111111";
                when x"D51" => data <= "1111111111";
                when x"D52" => data <= "1111111111";
                when x"D53" => data <= "1111111111";
                when x"D54" => data <= "1111111111";
                when x"D55" => data <= "1111111111";
                when x"D56" => data <= "1111111111";
                when x"D57" => data <= "1111111111";
                when x"D58" => data <= "1111111111";
                when x"D59" => data <= "1111111111";
                when x"D5A" => data <= "1111111111";
                when x"D5B" => data <= "1111111111";
                when x"D5C" => data <= "1111111111";
                when x"D5D" => data <= "1111111111";
                when x"D5E" => data <= "1111111111";
                when x"D5F" => data <= "1111111111";
                when x"D60" => data <= "1111111111";
                when x"D61" => data <= "1111111111";
                when x"D62" => data <= "1111111111";
                when x"D63" => data <= "1111111111";
                when x"D64" => data <= "1111111111";
                when x"D65" => data <= "1111111111";
                when x"D66" => data <= "1111111111";
                when x"D67" => data <= "1111111111";
                when x"D68" => data <= "1111111111";
                when x"D69" => data <= "1111111111";
                when x"D6A" => data <= "1111111111";
                when x"D6B" => data <= "1111111111";
                when x"D6C" => data <= "1111111111";
                when x"D6D" => data <= "1111111111";
                when x"D6E" => data <= "1111111111";
                when x"D6F" => data <= "1111111111";
                when x"D70" => data <= "1111111111";
                when x"D71" => data <= "1111111111";
                when x"D72" => data <= "1111111111";
                when x"D73" => data <= "1111111111";
                when x"D74" => data <= "1111111111";
                when x"D75" => data <= "1111111111";
                when x"D76" => data <= "1111111111";
                when x"D77" => data <= "1111111111";
                when x"D78" => data <= "1111111111";
                when x"D79" => data <= "1111111111";
                when x"D7A" => data <= "1111111111";
                when x"D7B" => data <= "1111111111";
                when x"D7C" => data <= "1111111111";
                when x"D7D" => data <= "1111111111";
                when x"D7E" => data <= "1111111111";
                when x"D7F" => data <= "1111111111";
                when x"D80" => data <= "1111111111";
                when x"D81" => data <= "1111111111";
                when x"D82" => data <= "1111111111";
                when x"D83" => data <= "1111111111";
                when x"D84" => data <= "1111111111";
                when x"D85" => data <= "1111111111";
                when x"D86" => data <= "1111111111";
                when x"D87" => data <= "1111111111";
                when x"D88" => data <= "1111111111";
                when x"D89" => data <= "1111111111";
                when x"D8A" => data <= "1111111111";
                when x"D8B" => data <= "1111111111";
                when x"D8C" => data <= "1111111111";
                when x"D8D" => data <= "1111111111";
                when x"D8E" => data <= "1111111111";
                when x"D8F" => data <= "1111111111";
                when x"D90" => data <= "1111111111";
                when x"D91" => data <= "1111111111";
                when x"D92" => data <= "1111111111";
                when x"D93" => data <= "1111111111";
                when x"D94" => data <= "1111111111";
                when x"D95" => data <= "1111111111";
                when x"D96" => data <= "1111111111";
                when x"D97" => data <= "1111111111";
                when x"D98" => data <= "1111111111";
                when x"D99" => data <= "1111111111";
                when x"D9A" => data <= "1111111111";
                when x"D9B" => data <= "1111111111";
                when x"D9C" => data <= "1111111111";
                when x"D9D" => data <= "1111111111";
                when x"D9E" => data <= "1111111111";
                when x"D9F" => data <= "1111111111";
                when x"DA0" => data <= "1111111111";
                when x"DA1" => data <= "1111111111";
                when x"DA2" => data <= "1111111111";
                when x"DA3" => data <= "1111111111";
                when x"DA4" => data <= "1111111111";
                when x"DA5" => data <= "1111111111";
                when x"DA6" => data <= "1111111111";
                when x"DA7" => data <= "1111111111";
                when x"DA8" => data <= "1111111111";
                when x"DA9" => data <= "1111111111";
                when x"DAA" => data <= "1111111111";
                when x"DAB" => data <= "1111111111";
                when x"DAC" => data <= "1111111111";
                when x"DAD" => data <= "1111111111";
                when x"DAE" => data <= "1111111111";
                when x"DAF" => data <= "1111111111";
                when x"DB0" => data <= "1111111111";
                when x"DB1" => data <= "1111111111";
                when x"DB2" => data <= "1111111111";
                when x"DB3" => data <= "1111111111";
                when x"DB4" => data <= "1111111111";
                when x"DB5" => data <= "1111111111";
                when x"DB6" => data <= "1111111111";
                when x"DB7" => data <= "1111111111";
                when x"DB8" => data <= "1111111111";
                when x"DB9" => data <= "1111111111";
                when x"DBA" => data <= "1111111111";
                when x"DBB" => data <= "1111111111";
                when x"DBC" => data <= "1111111111";
                when x"DBD" => data <= "1111111111";
                when x"DBE" => data <= "1111111111";
                when x"DBF" => data <= "1111111111";
                when x"DC0" => data <= "1111111111";
                when x"DC1" => data <= "1111111111";
                when x"DC2" => data <= "1111111111";
                when x"DC3" => data <= "1111111111";
                when x"DC4" => data <= "1111111111";
                when x"DC5" => data <= "1111111111";
                when x"DC6" => data <= "1111111111";
                when x"DC7" => data <= "1111111111";
                when x"DC8" => data <= "1111111111";
                when x"DC9" => data <= "1111111111";
                when x"DCA" => data <= "1111111111";
                when x"DCB" => data <= "1111111111";
                when x"DCC" => data <= "1111111111";
                when x"DCD" => data <= "1111111111";
                when x"DCE" => data <= "1111111111";
                when x"DCF" => data <= "1111111111";
                when x"DD0" => data <= "1111111111";
                when x"DD1" => data <= "1111111111";
                when x"DD2" => data <= "1000001000";
                when x"DD3" => data <= "1111111111";
                when x"DD4" => data <= "1111111111";
                when x"DD5" => data <= "1111111111";
                when x"DD6" => data <= "1111111111";
                when x"DD7" => data <= "1111111111";
                when x"DD8" => data <= "1111111111";
                when x"DD9" => data <= "1111111111";
                when x"DDA" => data <= "1111111111";
                when x"DDB" => data <= "1111111111";
                when x"DDC" => data <= "1111111111";
                when x"DDD" => data <= "1111111111";
                when x"DDE" => data <= "1111111111";
                when x"DDF" => data <= "1111111111";
                when x"DE0" => data <= "1111111111";
                when x"DE1" => data <= "1111111111";
                when x"DE2" => data <= "1111111111";
                when x"DE3" => data <= "1000111101";
                when x"DE4" => data <= "1111111111";
                when x"DE5" => data <= "1111111111";
                when x"DE6" => data <= "1111111111";
                when x"DE7" => data <= "1111111111";
                when x"DE8" => data <= "1111111111";
                when x"DE9" => data <= "1111111111";
                when x"DEA" => data <= "1111111111";
                when x"DEB" => data <= "1111111111";
                when x"DEC" => data <= "1111111111";
                when x"DED" => data <= "1111111111";
                when x"DEE" => data <= "1111111111";
                when x"DEF" => data <= "1111111111";
                when x"DF0" => data <= "1111111111";
                when x"DF1" => data <= "1111111111";
                when x"DF2" => data <= "1111111111";
                when x"DF3" => data <= "1111111111";
                when x"DF4" => data <= "1111111111";
                when x"DF5" => data <= "1111111111";
                when x"DF6" => data <= "1111111111";
                when x"DF7" => data <= "1111111111";
                when x"DF8" => data <= "1111111111";
                when x"DF9" => data <= "1111111111";
                when x"DFA" => data <= "1111111111";
                when x"DFB" => data <= "1111111111";
                when x"DFC" => data <= "1111111111";
                when x"DFD" => data <= "1111111111";
                when x"DFE" => data <= "1111111111";
                when x"DFF" => data <= "1111111111";
                when x"E00" => data <= "1111111111";
                when x"E01" => data <= "1111111111";
                when x"E02" => data <= "1111111111";
                when x"E03" => data <= "1111111111";
                when x"E04" => data <= "1111111111";
                when x"E05" => data <= "1111111111";
                when x"E06" => data <= "1111111111";
                when x"E07" => data <= "1111111111";
                when x"E08" => data <= "1111111111";
                when x"E09" => data <= "1111111111";
                when x"E0A" => data <= "1111111111";
                when x"E0B" => data <= "1111111111";
                when x"E0C" => data <= "1111111111";
                when x"E0D" => data <= "1111111111";
                when x"E0E" => data <= "1111111111";
                when x"E0F" => data <= "1111111111";
                when x"E10" => data <= "1111111111";
                when x"E11" => data <= "1111111111";
                when x"E12" => data <= "1111111111";
                when x"E13" => data <= "1111111111";
                when x"E14" => data <= "1111111111";
                when x"E15" => data <= "1111111111";
                when x"E16" => data <= "1111111111";
                when x"E17" => data <= "1111111111";
                when x"E18" => data <= "1111111111";
                when x"E19" => data <= "1111111111";
                when x"E1A" => data <= "1111111111";
                when x"E1B" => data <= "1111111111";
                when x"E1C" => data <= "1111111111";
                when x"E1D" => data <= "1111111111";
                when x"E1E" => data <= "1111111111";
                when x"E1F" => data <= "1111111111";
                when x"E20" => data <= "1111111111";
                when x"E21" => data <= "0000100100";
                when x"E22" => data <= "1111111111";
                when x"E23" => data <= "1111111111";
                when x"E24" => data <= "1111111111";
                when x"E25" => data <= "1111111111";
                when x"E26" => data <= "1111111111";
                when x"E27" => data <= "1111111111";
                when x"E28" => data <= "1111111111";
                when x"E29" => data <= "1111111111";
                when x"E2A" => data <= "1111111111";
                when x"E2B" => data <= "1111111111";
                when x"E2C" => data <= "1111111111";
                when x"E2D" => data <= "1111111111";
                when x"E2E" => data <= "1111111111";
                when x"E2F" => data <= "1111111111";
                when x"E30" => data <= "1111111111";
                when x"E31" => data <= "1111111111";
                when x"E32" => data <= "1111111111";
                when x"E33" => data <= "1111111111";
                when x"E34" => data <= "1111111111";
                when x"E35" => data <= "1000001000";
                when x"E36" => data <= "1111111111";
                when x"E37" => data <= "1111111111";
                when x"E38" => data <= "1111111111";
                when x"E39" => data <= "1111111111";
                when x"E3A" => data <= "1111111111";
                when x"E3B" => data <= "1111111111";
                when x"E3C" => data <= "1111111111";
                when x"E3D" => data <= "1111111111";
                when x"E3E" => data <= "1111111111";
                when x"E3F" => data <= "1111111111";
                when x"E40" => data <= "1111111111";
                when x"E41" => data <= "1111111111";
                when x"E42" => data <= "1111111111";
                when x"E43" => data <= "1111111111";
                when x"E44" => data <= "1111111111";
                when x"E45" => data <= "1111111111";
                when x"E46" => data <= "1111111111";
                when x"E47" => data <= "1111111111";
                when x"E48" => data <= "1111111111";
                when x"E49" => data <= "1111111111";
                when x"E4A" => data <= "1111111111";
                when x"E4B" => data <= "1111111111";
                when x"E4C" => data <= "1111111111";
                when x"E4D" => data <= "1111111111";
                when x"E4E" => data <= "1111111111";
                when x"E4F" => data <= "1111111111";
                when x"E50" => data <= "1111111111";
                when x"E51" => data <= "1111111111";
                when x"E52" => data <= "1111111111";
                when x"E53" => data <= "1111111111";
                when x"E54" => data <= "1111111111";
                when x"E55" => data <= "1111111111";
                when x"E56" => data <= "1111111111";
                when x"E57" => data <= "1111111111";
                when x"E58" => data <= "1111111111";
                when x"E59" => data <= "1111111111";
                when x"E5A" => data <= "1111111111";
                when x"E5B" => data <= "1111111111";
                when x"E5C" => data <= "1111111111";
                when x"E5D" => data <= "1111111111";
                when x"E5E" => data <= "1111111111";
                when x"E5F" => data <= "1111111111";
                when x"E60" => data <= "1111111111";
                when x"E61" => data <= "1111111111";
                when x"E62" => data <= "1111111111";
                when x"E63" => data <= "1111111111";
                when x"E64" => data <= "1111111111";
                when x"E65" => data <= "1111111111";
                when x"E66" => data <= "1111111111";
                when x"E67" => data <= "1111111111";
                when x"E68" => data <= "1111111111";
                when x"E69" => data <= "1111111111";
                when x"E6A" => data <= "1111111111";
                when x"E6B" => data <= "1111111111";
                when x"E6C" => data <= "1111111111";
                when x"E6D" => data <= "1111111111";
                when x"E6E" => data <= "1111111111";
                when x"E6F" => data <= "1111111111";
                when x"E70" => data <= "1111111111";
                when x"E71" => data <= "1111111111";
                when x"E72" => data <= "1111111111";
                when x"E73" => data <= "1111111111";
                when x"E74" => data <= "1111111111";
                when x"E75" => data <= "1111111111";
                when x"E76" => data <= "1111111111";
                when x"E77" => data <= "1111111111";
                when x"E78" => data <= "1111111111";
                when x"E79" => data <= "1111111111";
                when x"E7A" => data <= "1111111111";
                when x"E7B" => data <= "0110001100";
                when x"E7C" => data <= "1111111111";
                when x"E7D" => data <= "1111111111";
                when x"E7E" => data <= "1111111111";
                when x"E7F" => data <= "1111111111";
                when x"E80" => data <= "1111111111";
                when x"E81" => data <= "1111111111";
                when x"E82" => data <= "1111111111";
                when x"E83" => data <= "1111111111";
                when x"E84" => data <= "1111111111";
                when x"E85" => data <= "1111111111";
                when x"E86" => data <= "1111111111";
                when x"E87" => data <= "1111111111";
                when x"E88" => data <= "1111111111";
                when x"E89" => data <= "1111111111";
                when x"E8A" => data <= "1111111111";
                when x"E8B" => data <= "1111111111";
                when x"E8C" => data <= "1111111111";
                when x"E8D" => data <= "1111111111";
                when x"E8E" => data <= "1111111111";
                when x"E8F" => data <= "1111111111";
                when x"E90" => data <= "1111111111";
                when x"E91" => data <= "1111111111";
                when x"E92" => data <= "1111111111";
                when x"E93" => data <= "1111111111";
                when x"E94" => data <= "1111111111";
                when x"E95" => data <= "1111111111";
                when x"E96" => data <= "1111111111";
                when x"E97" => data <= "1111111111";
                when x"E98" => data <= "1111111111";
                when x"E99" => data <= "1111111111";
                when x"E9A" => data <= "1111111111";
                when x"E9B" => data <= "1111111111";
                when x"E9C" => data <= "1111111111";
                when x"E9D" => data <= "1111111111";
                when x"E9E" => data <= "1111111111";
                when x"E9F" => data <= "1111111111";
                when x"EA0" => data <= "1111111111";
                when x"EA1" => data <= "1111111111";
                when x"EA2" => data <= "1111111111";
                when x"EA3" => data <= "1111111111";
                when x"EA4" => data <= "1111111111";
                when x"EA5" => data <= "1111111111";
                when x"EA6" => data <= "1111111111";
                when x"EA7" => data <= "1111111111";
                when x"EA8" => data <= "1111111111";
                when x"EA9" => data <= "1111111111";
                when x"EAA" => data <= "1111111111";
                when x"EAB" => data <= "1111111111";
                when x"EAC" => data <= "1111111111";
                when x"EAD" => data <= "1111111111";
                when x"EAE" => data <= "1111111111";
                when x"EAF" => data <= "1111111111";
                when x"EB0" => data <= "1111111111";
                when x"EB1" => data <= "1111111111";
                when x"EB2" => data <= "1111111111";
                when x"EB3" => data <= "1111111111";
                when x"EB4" => data <= "1111111111";
                when x"EB5" => data <= "1000001000";
                when x"EB6" => data <= "1111111111";
                when x"EB7" => data <= "1111111111";
                when x"EB8" => data <= "1111111111";
                when x"EB9" => data <= "1111111111";
                when x"EBA" => data <= "1111111111";
                when x"EBB" => data <= "1111111111";
                when x"EBC" => data <= "1111111111";
                when x"EBD" => data <= "1111111111";
                when x"EBE" => data <= "1111111111";
                when x"EBF" => data <= "1111111111";
                when x"EC0" => data <= "1111111111";
                when x"EC1" => data <= "1111111111";
                when x"EC2" => data <= "1111111111";
                when x"EC3" => data <= "1111111111";
                when x"EC4" => data <= "1111111111";
                when x"EC5" => data <= "1111111111";
                when x"EC6" => data <= "1111111111";
                when x"EC7" => data <= "1111111111";
                when x"EC8" => data <= "1111111111";
                when x"EC9" => data <= "1111111111";
                when x"ECA" => data <= "1111111111";
                when x"ECB" => data <= "1111111111";
                when x"ECC" => data <= "1111111111";
                when x"ECD" => data <= "1111111111";
                when x"ECE" => data <= "1111111111";
                when x"ECF" => data <= "1111111111";
                when x"ED0" => data <= "1111111111";
                when x"ED1" => data <= "1111111111";
                when x"ED2" => data <= "1111111111";
                when x"ED3" => data <= "1111111111";
                when x"ED4" => data <= "1111111111";
                when x"ED5" => data <= "1111111111";
                when x"ED6" => data <= "1111111111";
                when x"ED7" => data <= "1111111111";
                when x"ED8" => data <= "1111111111";
                when x"ED9" => data <= "1111111111";
                when x"EDA" => data <= "1111111111";
                when x"EDB" => data <= "1111111111";
                when x"EDC" => data <= "1111111111";
                when x"EDD" => data <= "1111111111";
                when x"EDE" => data <= "1111111111";
                when x"EDF" => data <= "1111111111";
                when x"EE0" => data <= "1111111111";
                when x"EE1" => data <= "1111111111";
                when x"EE2" => data <= "1111111111";
                when x"EE3" => data <= "1111111111";
                when x"EE4" => data <= "1111111111";
                when x"EE5" => data <= "1111111111";
                when x"EE6" => data <= "1111111111";
                when x"EE7" => data <= "1111111111";
                when x"EE8" => data <= "1111111111";
                when x"EE9" => data <= "1111111111";
                when x"EEA" => data <= "1111111111";
                when x"EEB" => data <= "1111111111";
                when x"EEC" => data <= "1111111111";
                when x"EED" => data <= "1111111111";
                when x"EEE" => data <= "1111111111";
                when x"EEF" => data <= "1111111111";
                when x"EF0" => data <= "1111111111";
                when x"EF1" => data <= "1111111111";
                when x"EF2" => data <= "1111111111";
                when x"EF3" => data <= "1111111111";
                when x"EF4" => data <= "1111111111";
                when x"EF5" => data <= "1111111111";
                when x"EF6" => data <= "1111111111";
                when x"EF7" => data <= "1111111111";
                when x"EF8" => data <= "1111111111";
                when x"EF9" => data <= "1111111111";
                when x"EFA" => data <= "1111111111";
                when x"EFB" => data <= "1111111111";
                when x"EFC" => data <= "1111111111";
                when x"EFD" => data <= "1111111111";
                when x"EFE" => data <= "1111111111";
                when x"EFF" => data <= "1111111111";
                when x"F00" => data <= "1111111111";
                when x"F01" => data <= "1111111111";
                when x"F02" => data <= "1111111111";
                when x"F03" => data <= "1111111111";
                when x"F04" => data <= "1111111111";
                when x"F05" => data <= "1111111111";
                when x"F06" => data <= "1111111111";
                when x"F07" => data <= "1111111111";
                when x"F08" => data <= "1111111111";
                when x"F09" => data <= "1000001000";
                when x"F0A" => data <= "1111111111";
                when x"F0B" => data <= "1111111111";
                when x"F0C" => data <= "1111111111";
                when x"F0D" => data <= "1111111111";
                when x"F0E" => data <= "1111111111";
                when x"F0F" => data <= "1111111111";
                when x"F10" => data <= "1111111111";
                when x"F11" => data <= "1111111111";
                when x"F12" => data <= "1111111111";
                when x"F13" => data <= "1111111111";
                when x"F14" => data <= "1111111111";
                when x"F15" => data <= "1111111111";
                when x"F16" => data <= "1111111111";
                when x"F17" => data <= "1111111111";
                when x"F18" => data <= "1111111111";
                when x"F19" => data <= "1111111111";
                when x"F1A" => data <= "1111111111";
                when x"F1B" => data <= "1111111111";
                when x"F1C" => data <= "1111111111";
                when x"F1D" => data <= "1111111111";
                when x"F1E" => data <= "1111111111";
                when x"F1F" => data <= "1111111111";
                when x"F20" => data <= "1111111111";
                when x"F21" => data <= "1111111111";
                when x"F22" => data <= "1111111111";
                when x"F23" => data <= "1111111111";
                when x"F24" => data <= "1111111111";
                when x"F25" => data <= "1111111111";
                when x"F26" => data <= "1111111111";
                when x"F27" => data <= "1111111111";
                when x"F28" => data <= "1111111111";
                when x"F29" => data <= "1111111111";
                when x"F2A" => data <= "1111111111";
                when x"F2B" => data <= "1111111111";
                when x"F2C" => data <= "1111111111";
                when x"F2D" => data <= "1111111111";
                when x"F2E" => data <= "1111111111";
                when x"F2F" => data <= "1111111111";
                when x"F30" => data <= "1111111111";
                when x"F31" => data <= "1111111111";
                when x"F32" => data <= "1111111111";
                when x"F33" => data <= "1111111111";
                when x"F34" => data <= "1000001000";
                when x"F35" => data <= "1111111111";
                when x"F36" => data <= "1111111111";
                when x"F37" => data <= "1111111111";
                when x"F38" => data <= "1111111111";
                when x"F39" => data <= "1111111111";
                when x"F3A" => data <= "1111111111";
                when x"F3B" => data <= "1111111111";
                when x"F3C" => data <= "1111111111";
                when x"F3D" => data <= "1111111111";
                when x"F3E" => data <= "1111111111";
                when x"F3F" => data <= "1111111111";
                when x"F40" => data <= "1111111111";
                when x"F41" => data <= "1111111111";
                when x"F42" => data <= "1111111111";
                when x"F43" => data <= "1111111111";
                when x"F44" => data <= "1111111111";
                when x"F45" => data <= "1111111111";
                when x"F46" => data <= "1111111111";
                when x"F47" => data <= "1111111111";
                when x"F48" => data <= "1111111111";
                when x"F49" => data <= "1111111111";
                when x"F4A" => data <= "1111111111";
                when x"F4B" => data <= "1111111111";
                when x"F4C" => data <= "1111111111";
                when x"F4D" => data <= "1111111111";
                when x"F4E" => data <= "1111111111";
                when x"F4F" => data <= "1111111111";
                when x"F50" => data <= "1111111111";
                when x"F51" => data <= "1111111111";
                when x"F52" => data <= "1111111111";
                when x"F53" => data <= "1111111111";
                when x"F54" => data <= "1111111111";
                when x"F55" => data <= "1111111111";
                when x"F56" => data <= "1111111111";
                when x"F57" => data <= "1111111111";
                when x"F58" => data <= "1111111111";
                when x"F59" => data <= "1111111111";
                when x"F5A" => data <= "1111111111";
                when x"F5B" => data <= "1111111111";
                when x"F5C" => data <= "1111111111";
                when x"F5D" => data <= "1111111111";
                when x"F5E" => data <= "1111111111";
                when x"F5F" => data <= "1111111111";
                when x"F60" => data <= "1111111111";
                when x"F61" => data <= "1111111111";
                when x"F62" => data <= "1000001000";
                when x"F63" => data <= "1111111111";
                when x"F64" => data <= "1111111111";
                when x"F65" => data <= "1111111111";
                when x"F66" => data <= "1111111111";
                when x"F67" => data <= "1111111111";
                when x"F68" => data <= "1111111111";
                when x"F69" => data <= "1111111111";
                when x"F6A" => data <= "1111111111";
                when x"F6B" => data <= "1111111111";
                when x"F6C" => data <= "1111111111";
                when x"F6D" => data <= "1111111111";
                when x"F6E" => data <= "1111111111";
                when x"F6F" => data <= "1111111111";
                when x"F70" => data <= "1111111111";
                when x"F71" => data <= "1111111111";
                when x"F72" => data <= "1111111111";
                when x"F73" => data <= "1111111111";
                when x"F74" => data <= "1111111111";
                when x"F75" => data <= "1111111111";
                when x"F76" => data <= "1111111111";
                when x"F77" => data <= "1111111111";
                when x"F78" => data <= "1111111111";
                when x"F79" => data <= "1111111111";
                when x"F7A" => data <= "1111111111";
                when x"F7B" => data <= "1111111111";
                when x"F7C" => data <= "1111111111";
                when x"F7D" => data <= "1111111111";
                when x"F7E" => data <= "1111111111";
                when x"F7F" => data <= "1111111111";
                when x"F80" => data <= "1111111111";
                when x"F81" => data <= "1111111111";
                when x"F82" => data <= "1111111111";
                when x"F83" => data <= "1111111111";
                when x"F84" => data <= "1111111111";
                when x"F85" => data <= "1111111111";
                when x"F86" => data <= "1111111111";
                when x"F87" => data <= "1111111111";
                when x"F88" => data <= "1111111111";
                when x"F89" => data <= "1111111111";
                when x"F8A" => data <= "1111111111";
                when x"F8B" => data <= "1111111111";
                when x"F8C" => data <= "1111111111";
                when x"F8D" => data <= "1111111111";
                when x"F8E" => data <= "1111111111";
                when x"F8F" => data <= "1111111111";
                when x"F90" => data <= "1111111111";
                when x"F91" => data <= "1111111111";
                when x"F92" => data <= "1111111111";
                when x"F93" => data <= "1111111111";
                when x"F94" => data <= "1111111111";
                when x"F95" => data <= "1111111111";
                when x"F96" => data <= "1111111111";
                when x"F97" => data <= "1111111111";
                when x"F98" => data <= "1111111111";
                when x"F99" => data <= "1111111111";
                when x"F9A" => data <= "1111111111";
                when x"F9B" => data <= "1111111111";
                when x"F9C" => data <= "1111111111";
                when x"F9D" => data <= "1111111111";
                when x"F9E" => data <= "1111111111";
                when x"F9F" => data <= "1111111111";
                when x"FA0" => data <= "1111111111";
                when x"FA1" => data <= "1111111111";
                when x"FA2" => data <= "1111111111";
                when x"FA3" => data <= "1111111111";
                when x"FA4" => data <= "1111111111";
                when x"FA5" => data <= "1111111111";
                when x"FA6" => data <= "1111111111";
                when x"FA7" => data <= "1111111111";
                when x"FA8" => data <= "1111111111";
                when x"FA9" => data <= "1111111111";
                when x"FAA" => data <= "1111111111";
                when x"FAB" => data <= "1111111111";
                when x"FAC" => data <= "1111111111";
                when x"FAD" => data <= "1111111111";
                when x"FAE" => data <= "1111111111";
                when x"FAF" => data <= "1111111111";
                when x"FB0" => data <= "1111111111";
                when x"FB1" => data <= "1111111111";
                when x"FB2" => data <= "1111111111";
                when x"FB3" => data <= "1111111111";
                when x"FB4" => data <= "1111111111";
                when x"FB5" => data <= "1111111111";
                when x"FB6" => data <= "1111111111";
                when x"FB7" => data <= "1111111111";
                when x"FB8" => data <= "1111111111";
                when x"FB9" => data <= "1111111111";
                when x"FBA" => data <= "0100000111";
                when x"FBB" => data <= "1111111111";
                when x"FBC" => data <= "1111111111";
                when x"FBD" => data <= "1111111111";
                when x"FBE" => data <= "1000001000";
                when x"FBF" => data <= "1111111111";
                when x"FC0" => data <= "1111111111";
                when x"FC1" => data <= "1111111111";
                when x"FC2" => data <= "1111111111";
                when x"FC3" => data <= "1111111111";
                when x"FC4" => data <= "1111111111";
                when x"FC5" => data <= "1111111111";
                when x"FC6" => data <= "1111111111";
                when x"FC7" => data <= "1111111111";
                when x"FC8" => data <= "1111111111";
                when x"FC9" => data <= "1111111111";
                when x"FCA" => data <= "1111111111";
                when x"FCB" => data <= "1111111111";
                when x"FCC" => data <= "1111111111";
                when x"FCD" => data <= "1111111111";
                when x"FCE" => data <= "1111111111";
                when x"FCF" => data <= "1111111111";
                when x"FD0" => data <= "1111111111";
                when x"FD1" => data <= "1111111111";
                when x"FD2" => data <= "1111111111";
                when x"FD3" => data <= "1111111111";
                when x"FD4" => data <= "1111111111";
                when x"FD5" => data <= "1111111111";
                when x"FD6" => data <= "1111111111";
                when x"FD7" => data <= "1111111111";
                when x"FD8" => data <= "1111111111";
                when x"FD9" => data <= "1111111111";
                when x"FDA" => data <= "1111111111";
                when x"FDB" => data <= "1111111111";
                when x"FDC" => data <= "1111111111";
                when x"FDD" => data <= "1111111111";
                when x"FDE" => data <= "1111111111";
                when x"FDF" => data <= "1111111111";
                when x"FE0" => data <= "1111111111";
                when x"FE1" => data <= "1111111111";
                when x"FE2" => data <= "1111111111";
                when x"FE3" => data <= "1111111111";
                when x"FE4" => data <= "1111111111";
                when x"FE5" => data <= "1111111111";
                when x"FE6" => data <= "1111111111";
                when x"FE7" => data <= "1111111111";
                when x"FE8" => data <= "1111111111";
                when x"FE9" => data <= "1111111111";
                when x"FEA" => data <= "1111111111";
                when x"FEB" => data <= "1111111111";
                when x"FEC" => data <= "1111111111";
                when x"FED" => data <= "1111111111";
                when x"FEE" => data <= "1111111111";
                when x"FEF" => data <= "1111111111";
                when x"FF0" => data <= "1111111111";
                when x"FF1" => data <= "1111111111";
                when x"FF2" => data <= "1111111111";
                when x"FF3" => data <= "1111111111";
                when x"FF4" => data <= "1111111111";
                when x"FF5" => data <= "1111111111";
                when x"FF6" => data <= "1111111111";
                when x"FF7" => data <= "1111111111";
                when x"FF8" => data <= "1111111111";
                when x"FF9" => data <= "1111111111";
                when x"FFA" => data <= "1111111111";
                when x"FFB" => data <= "1111111111";
                when x"FFC" => data <= "1111111111";
                when x"FFD" => data <= "1111111111";
                when x"FFE" => data <= "1111111111";
                when x"FFF" => data <= "1111111111";
                when x"1000" => data <= "1111111111";
                when x"1001" => data <= "1111111111";
                when x"1002" => data <= "1111111111";
                when x"1003" => data <= "1111111111";
                when x"1004" => data <= "1111111111";
                when x"1005" => data <= "1111111111";
                when x"1006" => data <= "1111111111";
                when x"1007" => data <= "1111111111";
                when x"1008" => data <= "1111111111";
                when x"1009" => data <= "1111111111";
                when x"100A" => data <= "1111111111";
                when x"100B" => data <= "1111111111";
                when x"100C" => data <= "1111111111";
                when x"100D" => data <= "1111111111";
                when x"100E" => data <= "1111111111";
                when x"100F" => data <= "1111111111";
                when x"1010" => data <= "1111111111";
                when x"1011" => data <= "1111111111";
                when x"1012" => data <= "1111111111";
                when x"1013" => data <= "1111111111";
                when x"1014" => data <= "1111111111";
                when x"1015" => data <= "1111111111";
                when x"1016" => data <= "1111111111";
                when x"1017" => data <= "1111111111";
                when x"1018" => data <= "1111111111";
                when x"1019" => data <= "1111111111";
                when x"101A" => data <= "1111111111";
                when x"101B" => data <= "1111111111";
                when x"101C" => data <= "1111111111";
                when x"101D" => data <= "1111111111";
                when x"101E" => data <= "1111111111";
                when x"101F" => data <= "1111111111";
                when x"1020" => data <= "1111111111";
                when x"1021" => data <= "1111111111";
                when x"1022" => data <= "1111111111";
                when x"1023" => data <= "1111111111";
                when x"1024" => data <= "1111111111";
                when x"1025" => data <= "1111111111";
                when x"1026" => data <= "1111111111";
                when x"1027" => data <= "1111111111";
                when x"1028" => data <= "1111111111";
                when x"1029" => data <= "1111111111";
                when x"102A" => data <= "1111111111";
                when x"102B" => data <= "1111111111";
                when x"102C" => data <= "1111111111";
                when x"102D" => data <= "1111111111";
                when x"102E" => data <= "1111111111";
                when x"102F" => data <= "1111111111";
                when x"1030" => data <= "1111111111";
                when x"1031" => data <= "1111111111";
                when x"1032" => data <= "1111111111";
                when x"1033" => data <= "1111111111";
                when x"1034" => data <= "1111111111";
                when x"1035" => data <= "1111111111";
                when x"1036" => data <= "1111111111";
                when x"1037" => data <= "1111111111";
                when x"1038" => data <= "1111111111";
                when x"1039" => data <= "1111111111";
                when x"103A" => data <= "1111111111";
                when x"103B" => data <= "1111111111";
                when x"103C" => data <= "1111111111";
                when x"103D" => data <= "1111111111";
                when x"103E" => data <= "1111111111";
                when x"103F" => data <= "1111111111";
                when x"1040" => data <= "1111111111";
                when x"1041" => data <= "1111111111";
                when x"1042" => data <= "1111111111";
                when x"1043" => data <= "1111111111";
                when x"1044" => data <= "1111111111";
                when x"1045" => data <= "1111111111";
                when x"1046" => data <= "1111111111";
                when x"1047" => data <= "1111111111";
                when x"1048" => data <= "1111111111";
                when x"1049" => data <= "1111111111";
                when x"104A" => data <= "1111111111";
                when x"104B" => data <= "1111111111";
                when x"104C" => data <= "1111111111";
                when x"104D" => data <= "1111111111";
                when x"104E" => data <= "1111111111";
                when x"104F" => data <= "1111111111";
                when x"1050" => data <= "1111111111";
                when x"1051" => data <= "1111111111";
                when x"1052" => data <= "1111111111";
                when x"1053" => data <= "1111111111";
                when x"1054" => data <= "1111111111";
                when x"1055" => data <= "1111111111";
                when x"1056" => data <= "1111111111";
                when x"1057" => data <= "1111111111";
                when x"1058" => data <= "1111111111";
                when x"1059" => data <= "1111111111";
                when x"105A" => data <= "1111111111";
                when x"105B" => data <= "1111111111";
                when x"105C" => data <= "1111111111";
                when x"105D" => data <= "1111111111";
                when x"105E" => data <= "1111111111";
                when x"105F" => data <= "1111111111";
                when x"1060" => data <= "1111111111";
                when x"1061" => data <= "1111111111";
                when x"1062" => data <= "1111111111";
                when x"1063" => data <= "1111111111";
                when x"1064" => data <= "1111111111";
                when x"1065" => data <= "1111111111";
                when x"1066" => data <= "1111111111";
                when x"1067" => data <= "1111111111";
                when x"1068" => data <= "1111111111";
                when x"1069" => data <= "1111111111";
                when x"106A" => data <= "1111111111";
                when x"106B" => data <= "1111111111";
                when x"106C" => data <= "1111111111";
                when x"106D" => data <= "1111111111";
                when x"106E" => data <= "1111111111";
                when x"106F" => data <= "1111111111";
                when x"1070" => data <= "1111111111";
                when x"1071" => data <= "1111111111";
                when x"1072" => data <= "1111111111";
                when x"1073" => data <= "1111111111";
                when x"1074" => data <= "1111111111";
                when x"1075" => data <= "1111111111";
                when x"1076" => data <= "1111111111";
                when x"1077" => data <= "1111111111";
                when x"1078" => data <= "1111111111";
                when x"1079" => data <= "1111111111";
                when x"107A" => data <= "1111111111";
                when x"107B" => data <= "1111111111";
                when x"107C" => data <= "1111111111";
                when x"107D" => data <= "1111111111";
                when x"107E" => data <= "1111111111";
                when x"107F" => data <= "1111111111";
                when x"1080" => data <= "1111111111";
                when x"1081" => data <= "1111111111";
                when x"1082" => data <= "1111111111";
                when x"1083" => data <= "1111111111";
                when x"1084" => data <= "1111111111";
                when x"1085" => data <= "1111111111";
                when x"1086" => data <= "1111111111";
                when x"1087" => data <= "1111111111";
                when x"1088" => data <= "1111111111";
                when x"1089" => data <= "1111111111";
                when x"108A" => data <= "1111111111";
                when x"108B" => data <= "1111111111";
                when x"108C" => data <= "1111111111";
                when x"108D" => data <= "1111111111";
                when x"108E" => data <= "1111111111";
                when x"108F" => data <= "1111111111";
                when x"1090" => data <= "1111111111";
                when x"1091" => data <= "1000001000";
                when x"1092" => data <= "1111111111";
                when x"1093" => data <= "1111111111";
                when x"1094" => data <= "1111111111";
                when x"1095" => data <= "1111111111";
                when x"1096" => data <= "1111111111";
                when x"1097" => data <= "1111111111";
                when x"1098" => data <= "1000001000";
                when x"1099" => data <= "1111111111";
                when x"109A" => data <= "1111111111";
                when x"109B" => data <= "1111111111";
                when x"109C" => data <= "1111111111";
                when x"109D" => data <= "1111111111";
                when x"109E" => data <= "1111111111";
                when x"109F" => data <= "1111111111";
                when x"10A0" => data <= "1111111111";
                when x"10A1" => data <= "1111111111";
                when x"10A2" => data <= "1111111111";
                when x"10A3" => data <= "1111111111";
                when x"10A4" => data <= "1111111111";
                when x"10A5" => data <= "1111111111";
                when x"10A6" => data <= "1111111111";
                when x"10A7" => data <= "1111111111";
                when x"10A8" => data <= "1111111111";
                when x"10A9" => data <= "1111111111";
                when x"10AA" => data <= "1111111111";
                when x"10AB" => data <= "1011011100";
                when x"10AC" => data <= "1111111111";
                when x"10AD" => data <= "1111111111";
                when x"10AE" => data <= "1111111111";
                when x"10AF" => data <= "1111111111";
                when x"10B0" => data <= "1111111111";
                when x"10B1" => data <= "1111111111";
                when x"10B2" => data <= "1111111111";
                when x"10B3" => data <= "1111111111";
                when x"10B4" => data <= "1111111111";
                when x"10B5" => data <= "1111111111";
                when x"10B6" => data <= "1111111111";
                when x"10B7" => data <= "1111111111";
                when x"10B8" => data <= "1111111111";
                when x"10B9" => data <= "1111111111";
                when x"10BA" => data <= "1111111111";
                when x"10BB" => data <= "1111111111";
                when x"10BC" => data <= "1111111111";
                when x"10BD" => data <= "1111111111";
                when x"10BE" => data <= "1111111111";
                when x"10BF" => data <= "1111111111";
                when x"10C0" => data <= "1111111111";
                when x"10C1" => data <= "1111111111";
                when x"10C2" => data <= "1111111111";
                when x"10C3" => data <= "1111111111";
                when x"10C4" => data <= "1111111111";
                when x"10C5" => data <= "1111111111";
                when x"10C6" => data <= "1111111111";
                when x"10C7" => data <= "1111111111";
                when x"10C8" => data <= "1111111111";
                when x"10C9" => data <= "1111111111";
                when x"10CA" => data <= "1111111111";
                when x"10CB" => data <= "1111111111";
                when x"10CC" => data <= "1111111111";
                when x"10CD" => data <= "1111111111";
                when x"10CE" => data <= "0000100100";
                when x"10CF" => data <= "1111111111";
                when x"10D0" => data <= "0010101111";
                when x"10D1" => data <= "1111111111";
                when x"10D2" => data <= "1111111111";
                when x"10D3" => data <= "1111111111";
                when x"10D4" => data <= "1111111111";
                when x"10D5" => data <= "1111111111";
                when x"10D6" => data <= "1111111111";
                when x"10D7" => data <= "1111111111";
                when x"10D8" => data <= "1111111111";
                when x"10D9" => data <= "1111111111";
                when x"10DA" => data <= "1111111111";
                when x"10DB" => data <= "1111111111";
                when x"10DC" => data <= "1111111111";
                when x"10DD" => data <= "1111111111";
                when x"10DE" => data <= "1111111111";
                when x"10DF" => data <= "1111111111";
                when x"10E0" => data <= "1111111111";
                when x"10E1" => data <= "1111111111";
                when x"10E2" => data <= "1111111111";
                when x"10E3" => data <= "1111111111";
                when x"10E4" => data <= "1111111111";
                when x"10E5" => data <= "1111111111";
                when x"10E6" => data <= "1111111111";
                when x"10E7" => data <= "1111111111";
                when x"10E8" => data <= "1111111111";
                when x"10E9" => data <= "1111111111";
                when x"10EA" => data <= "1111111111";
                when x"10EB" => data <= "1111111111";
                when x"10EC" => data <= "1111111111";
                when x"10ED" => data <= "1111111111";
                when x"10EE" => data <= "1111111111";
                when x"10EF" => data <= "1111111111";
                when x"10F0" => data <= "1111111111";
                when x"10F1" => data <= "1111111111";
                when x"10F2" => data <= "1111111111";
                when x"10F3" => data <= "1111111111";
                when x"10F4" => data <= "1111111111";
                when x"10F5" => data <= "1111111111";
                when x"10F6" => data <= "1111111111";
                when x"10F7" => data <= "1111111111";
                when x"10F8" => data <= "1111111111";
                when x"10F9" => data <= "1111111111";
                when x"10FA" => data <= "1111111111";
                when x"10FB" => data <= "1111111111";
                when x"10FC" => data <= "1111111111";
                when x"10FD" => data <= "1111111111";
                when x"10FE" => data <= "1111111111";
                when x"10FF" => data <= "1111111111";
                when x"1100" => data <= "1111111111";
                when x"1101" => data <= "1111111111";
                when x"1102" => data <= "1111111111";
                when x"1103" => data <= "1111111111";
                when x"1104" => data <= "1111111111";
                when x"1105" => data <= "1111111111";
                when x"1106" => data <= "1111111111";
                when x"1107" => data <= "1111111111";
                when x"1108" => data <= "1111111111";
                when x"1109" => data <= "1111111111";
                when x"110A" => data <= "0000100100";
                when x"110B" => data <= "1111111111";
                when x"110C" => data <= "1111111111";
                when x"110D" => data <= "1111111111";
                when x"110E" => data <= "1111111111";
                when x"110F" => data <= "1111111111";
                when x"1110" => data <= "1111111111";
                when x"1111" => data <= "1111111111";
                when x"1112" => data <= "1111111111";
                when x"1113" => data <= "1111111111";
                when x"1114" => data <= "1111111111";
                when x"1115" => data <= "1111111111";
                when x"1116" => data <= "1111111111";
                when x"1117" => data <= "1111111111";
                when x"1118" => data <= "1111111111";
                when x"1119" => data <= "1111111111";
                when x"111A" => data <= "1111111111";
                when x"111B" => data <= "1111111111";
                when x"111C" => data <= "1111111111";
                when x"111D" => data <= "1111111111";
                when x"111E" => data <= "1111111111";
                when x"111F" => data <= "1111111111";
                when x"1120" => data <= "1111111111";
                when x"1121" => data <= "1111111111";
                when x"1122" => data <= "1111111111";
                when x"1123" => data <= "1111111111";
                when x"1124" => data <= "1111111111";
                when x"1125" => data <= "1111111111";
                when x"1126" => data <= "1111111111";
                when x"1127" => data <= "1111111111";
                when x"1128" => data <= "1111111111";
                when x"1129" => data <= "1111111111";
                when x"112A" => data <= "1111111111";
                when x"112B" => data <= "1111111111";
                when x"112C" => data <= "1111111111";
                when x"112D" => data <= "1111111111";
                when x"112E" => data <= "1111111111";
                when x"112F" => data <= "1111111111";
                when x"1130" => data <= "1111111111";
                when x"1131" => data <= "1111111111";
                when x"1132" => data <= "1111111111";
                when x"1133" => data <= "1111111111";
                when x"1134" => data <= "1111111111";
                when x"1135" => data <= "1111111111";
                when x"1136" => data <= "1111111111";
                when x"1137" => data <= "1111111111";
                when x"1138" => data <= "1111111111";
                when x"1139" => data <= "1111111111";
                when x"113A" => data <= "1111111111";
                when x"113B" => data <= "1111111111";
                when x"113C" => data <= "1111111111";
                when x"113D" => data <= "1111111111";
                when x"113E" => data <= "1111111111";
                when x"113F" => data <= "1111111111";
                when x"1140" => data <= "1111111111";
                when x"1141" => data <= "1111111111";
                when x"1142" => data <= "1111111111";
                when x"1143" => data <= "1111111111";
                when x"1144" => data <= "1111111111";
                when x"1145" => data <= "1111111111";
                when x"1146" => data <= "1111111111";
                when x"1147" => data <= "1111111111";
                when x"1148" => data <= "1111111111";
                when x"1149" => data <= "1111111111";
                when x"114A" => data <= "1111111111";
                when x"114B" => data <= "1111111111";
                when x"114C" => data <= "1111111111";
                when x"114D" => data <= "1111111111";
                when x"114E" => data <= "1111111111";
                when x"114F" => data <= "1111111111";
                when x"1150" => data <= "1111111111";
                when x"1151" => data <= "1111111111";
                when x"1152" => data <= "1111111111";
                when x"1153" => data <= "1111111111";
                when x"1154" => data <= "1111111111";
                when x"1155" => data <= "1000001000";
                when x"1156" => data <= "1111111111";
                when x"1157" => data <= "1111111111";
                when x"1158" => data <= "1111111111";
                when x"1159" => data <= "1111111111";
                when x"115A" => data <= "1111111111";
                when x"115B" => data <= "1111111111";
                when x"115C" => data <= "1111111111";
                when x"115D" => data <= "1111111111";
                when x"115E" => data <= "1111111111";
                when x"115F" => data <= "1111111111";
                when x"1160" => data <= "0001111011";
                when x"1161" => data <= "1111111111";
                when x"1162" => data <= "1111111111";
                when x"1163" => data <= "1111111111";
                when x"1164" => data <= "1111111111";
                when x"1165" => data <= "1111111111";
                when x"1166" => data <= "1111111111";
                when x"1167" => data <= "1111111111";
                when x"1168" => data <= "1111111111";
                when x"1169" => data <= "1111111111";
                when x"116A" => data <= "0100000111";
                when x"116B" => data <= "1111111111";
                when x"116C" => data <= "1111111111";
                when x"116D" => data <= "1111111111";
                when x"116E" => data <= "1111111111";
                when x"116F" => data <= "1111111111";
                when x"1170" => data <= "1111111111";
                when x"1171" => data <= "1111111111";
                when x"1172" => data <= "1111111111";
                when x"1173" => data <= "1111111111";
                when x"1174" => data <= "1111111111";
                when x"1175" => data <= "1111111111";
                when x"1176" => data <= "1111111111";
                when x"1177" => data <= "1111111111";
                when x"1178" => data <= "1111111111";
                when x"1179" => data <= "1111111111";
                when x"117A" => data <= "1111111111";
                when x"117B" => data <= "1111111111";
                when x"117C" => data <= "1111111111";
                when x"117D" => data <= "1111111111";
                when x"117E" => data <= "1111111111";
                when x"117F" => data <= "1111111111";
                when x"1180" => data <= "1111111111";
                when x"1181" => data <= "1111111111";
                when x"1182" => data <= "1111111111";
                when x"1183" => data <= "1111111111";
                when x"1184" => data <= "1111111111";
                when x"1185" => data <= "1111111111";
                when x"1186" => data <= "1111111111";
                when x"1187" => data <= "1111111111";
                when x"1188" => data <= "1111111111";
                when x"1189" => data <= "1111111111";
                when x"118A" => data <= "1111111111";
                when x"118B" => data <= "1111111111";
                when x"118C" => data <= "1111111111";
                when x"118D" => data <= "1111111111";
                when x"118E" => data <= "1111111111";
                when x"118F" => data <= "1111111111";
                when x"1190" => data <= "1111111111";
                when x"1191" => data <= "1111111111";
                when x"1192" => data <= "1111111111";
                when x"1193" => data <= "1111111111";
                when x"1194" => data <= "1111111111";
                when x"1195" => data <= "1111111111";
                when x"1196" => data <= "1111111111";
                when x"1197" => data <= "1111111111";
                when x"1198" => data <= "1111111111";
                when x"1199" => data <= "1111111111";
                when x"119A" => data <= "1111111111";
                when x"119B" => data <= "1111111111";
                when x"119C" => data <= "1111111111";
                when x"119D" => data <= "1111111111";
                when x"119E" => data <= "1111111111";
                when x"119F" => data <= "1111111111";
                when x"11A0" => data <= "1111111111";
                when x"11A1" => data <= "1111111111";
                when x"11A2" => data <= "1111111111";
                when x"11A3" => data <= "1111111111";
                when x"11A4" => data <= "1111111111";
                when x"11A5" => data <= "1111111111";
                when x"11A6" => data <= "1111111111";
                when x"11A7" => data <= "1111111111";
                when x"11A8" => data <= "1111111111";
                when x"11A9" => data <= "1111111111";
                when x"11AA" => data <= "1111111111";
                when x"11AB" => data <= "1111111111";
                when x"11AC" => data <= "1111111111";
                when x"11AD" => data <= "1111111111";
                when x"11AE" => data <= "1111111111";
                when x"11AF" => data <= "1111111111";
                when x"11B0" => data <= "1111111111";
                when x"11B1" => data <= "1111111111";
                when x"11B2" => data <= "1111111111";
                when x"11B3" => data <= "1111111111";
                when x"11B4" => data <= "1111111111";
                when x"11B5" => data <= "1111111111";
                when x"11B6" => data <= "1111111111";
                when x"11B7" => data <= "1111111111";
                when x"11B8" => data <= "1111111111";
                when x"11B9" => data <= "1111111111";
                when x"11BA" => data <= "1111111111";
                when x"11BB" => data <= "1111111111";
                when x"11BC" => data <= "1111111111";
                when x"11BD" => data <= "1111111111";
                when x"11BE" => data <= "1111111111";
                when x"11BF" => data <= "1111111111";
                when x"11C0" => data <= "1111111111";
                when x"11C1" => data <= "1111111111";
                when x"11C2" => data <= "1111111111";
                when x"11C3" => data <= "1111111111";
                when x"11C4" => data <= "1111111111";
                when x"11C5" => data <= "1111111111";
                when x"11C6" => data <= "1111111111";
                when x"11C7" => data <= "1111111111";
                when x"11C8" => data <= "1111111111";
                when x"11C9" => data <= "1111111111";
                when x"11CA" => data <= "1111111111";
                when x"11CB" => data <= "1111111111";
                when x"11CC" => data <= "1111111111";
                when x"11CD" => data <= "1111111111";
                when x"11CE" => data <= "1111111111";
                when x"11CF" => data <= "1111111111";
                when x"11D0" => data <= "1111111111";
                when x"11D1" => data <= "1111111111";
                when x"11D2" => data <= "1111111111";
                when x"11D3" => data <= "1111111111";
                when x"11D4" => data <= "1111111111";
                when x"11D5" => data <= "1111111111";
                when x"11D6" => data <= "1111111111";
                when x"11D7" => data <= "1111111111";
                when x"11D8" => data <= "1111111111";
                when x"11D9" => data <= "1111111111";
                when x"11DA" => data <= "1111111111";
                when x"11DB" => data <= "1111111111";
                when x"11DC" => data <= "1111111111";
                when x"11DD" => data <= "1111111111";
                when x"11DE" => data <= "1111111111";
                when x"11DF" => data <= "1111111111";
                when x"11E0" => data <= "1111111111";
                when x"11E1" => data <= "1111111111";
                when x"11E2" => data <= "1111111111";
                when x"11E3" => data <= "1111111111";
                when x"11E4" => data <= "1111111111";
                when x"11E5" => data <= "1111111111";
                when x"11E6" => data <= "1111111111";
                when x"11E7" => data <= "1111111111";
                when x"11E8" => data <= "1111111111";
                when x"11E9" => data <= "1111111111";
                when x"11EA" => data <= "1111111111";
                when x"11EB" => data <= "1111111111";
                when x"11EC" => data <= "1111111111";
                when x"11ED" => data <= "1111111111";
                when x"11EE" => data <= "1111111111";
                when x"11EF" => data <= "1111111111";
                when x"11F0" => data <= "1111111111";
                when x"11F1" => data <= "1111111111";
                when x"11F2" => data <= "1111111111";
                when x"11F3" => data <= "1111111111";
                when x"11F4" => data <= "1111111111";
                when x"11F5" => data <= "1111111111";
                when x"11F6" => data <= "1111111111";
                when x"11F7" => data <= "1111111111";
                when x"11F8" => data <= "1111111111";
                when x"11F9" => data <= "1111111111";
                when x"11FA" => data <= "1111111111";
                when x"11FB" => data <= "1111111111";
                when x"11FC" => data <= "1111111111";
                when x"11FD" => data <= "1111111111";
                when x"11FE" => data <= "1111111111";
                when x"11FF" => data <= "1111111111";
                when x"1200" => data <= "1111111111";
                when x"1201" => data <= "1111111111";
                when x"1202" => data <= "1111111111";
                when x"1203" => data <= "1111111111";
                when x"1204" => data <= "1111111111";
                when x"1205" => data <= "1111111111";
                when x"1206" => data <= "1111111111";
                when x"1207" => data <= "1111111111";
                when x"1208" => data <= "1111111111";
                when x"1209" => data <= "1111111111";
                when x"120A" => data <= "1111111111";
                when x"120B" => data <= "1111111111";
                when x"120C" => data <= "1111111111";
                when x"120D" => data <= "1111111111";
                when x"120E" => data <= "1111111111";
                when x"120F" => data <= "1111111111";
                when x"1210" => data <= "1111111111";
                when x"1211" => data <= "1111111111";
                when x"1212" => data <= "1000111101";
                when x"1213" => data <= "1111111111";
                when x"1214" => data <= "1111111111";
                when x"1215" => data <= "1111111111";
                when x"1216" => data <= "1111111111";
                when x"1217" => data <= "1111111111";
                when x"1218" => data <= "1111111111";
                when x"1219" => data <= "1111111111";
                when x"121A" => data <= "1111111111";
                when x"121B" => data <= "1111111111";
                when x"121C" => data <= "1111111111";
                when x"121D" => data <= "1111111111";
                when x"121E" => data <= "1111111111";
                when x"121F" => data <= "1111111111";
                when x"1220" => data <= "1111111111";
                when x"1221" => data <= "1111111111";
                when x"1222" => data <= "1111111111";
                when x"1223" => data <= "1111111111";
                when x"1224" => data <= "1111111111";
                when x"1225" => data <= "1111111111";
                when x"1226" => data <= "1111111111";
                when x"1227" => data <= "1111111111";
                when x"1228" => data <= "1111111111";
                when x"1229" => data <= "1111111111";
                when x"122A" => data <= "1111111111";
                when x"122B" => data <= "1111111111";
                when x"122C" => data <= "1111111111";
                when x"122D" => data <= "1111111111";
                when x"122E" => data <= "1111111111";
                when x"122F" => data <= "1111111111";
                when x"1230" => data <= "1111111111";
                when x"1231" => data <= "1111111111";
                when x"1232" => data <= "1111111111";
                when x"1233" => data <= "1111111111";
                when x"1234" => data <= "1111111111";
                when x"1235" => data <= "1111111111";
                when x"1236" => data <= "1111111111";
                when x"1237" => data <= "1111111111";
                when x"1238" => data <= "1111111111";
                when x"1239" => data <= "1111111111";
                when x"123A" => data <= "1111111111";
                when x"123B" => data <= "1111111111";
                when x"123C" => data <= "1111111111";
                when x"123D" => data <= "1111111111";
                when x"123E" => data <= "1111111111";
                when x"123F" => data <= "1111111111";
                when x"1240" => data <= "1111111111";
                when x"1241" => data <= "1111111111";
                when x"1242" => data <= "1111111111";
                when x"1243" => data <= "1111111111";
                when x"1244" => data <= "1111111111";
                when x"1245" => data <= "1111111111";
                when x"1246" => data <= "1111111111";
                when x"1247" => data <= "1111111111";
                when x"1248" => data <= "1111111111";
                when x"1249" => data <= "1111111111";
                when x"124A" => data <= "1111111111";
                when x"124B" => data <= "1111111111";
                when x"124C" => data <= "1111111111";
                when x"124D" => data <= "1111111111";
                when x"124E" => data <= "1111111111";
                when x"124F" => data <= "1111111111";
                when x"1250" => data <= "1111111111";
                when x"1251" => data <= "1111111111";
                when x"1252" => data <= "1111111111";
                when x"1253" => data <= "1000001000";
                when x"1254" => data <= "1111111111";
                when x"1255" => data <= "1111111111";
                when x"1256" => data <= "1111111111";
                when x"1257" => data <= "1111111111";
                when x"1258" => data <= "1111111111";
                when x"1259" => data <= "1111111111";
                when x"125A" => data <= "1111111111";
                when x"125B" => data <= "1111111111";
                when x"125C" => data <= "1111111111";
                when x"125D" => data <= "1111111111";
                when x"125E" => data <= "1111111111";
                when x"125F" => data <= "1111111111";
                when x"1260" => data <= "1111111111";
                when x"1261" => data <= "1111111111";
                when x"1262" => data <= "1111111111";
                when x"1263" => data <= "1111111111";
                when x"1264" => data <= "1111111111";
                when x"1265" => data <= "1111111111";
                when x"1266" => data <= "0010101111";
                when x"1267" => data <= "1111111111";
                when x"1268" => data <= "1111111111";
                when x"1269" => data <= "1111111111";
                when x"126A" => data <= "1111111111";
                when x"126B" => data <= "1111111111";
                when x"126C" => data <= "1111111111";
                when x"126D" => data <= "1111111111";
                when x"126E" => data <= "1111111111";
                when x"126F" => data <= "1111111111";
                when x"1270" => data <= "1111111111";
                when x"1271" => data <= "1111111111";
                when x"1272" => data <= "1111111111";
                when x"1273" => data <= "1111111111";
                when x"1274" => data <= "1111111111";
                when x"1275" => data <= "1111111111";
                when x"1276" => data <= "1111111111";
                when x"1277" => data <= "1111111111";
                when x"1278" => data <= "1111111111";
                when x"1279" => data <= "1111111111";
                when x"127A" => data <= "1111111111";
                when x"127B" => data <= "1111111111";
                when x"127C" => data <= "1111111111";
                when x"127D" => data <= "1111111111";
                when x"127E" => data <= "1111111111";
                when x"127F" => data <= "1111111111";
                when x"1280" => data <= "1111111111";
                when x"1281" => data <= "1111111111";
                when x"1282" => data <= "1111111111";
                when x"1283" => data <= "1111111111";
                when x"1284" => data <= "1111111111";
                when x"1285" => data <= "1111111111";
                when x"1286" => data <= "1111111111";
                when x"1287" => data <= "1111111111";
                when x"1288" => data <= "1111111111";
                when x"1289" => data <= "1111111111";
                when x"128A" => data <= "1111111111";
                when x"128B" => data <= "1111111111";
                when x"128C" => data <= "1111111111";
                when x"128D" => data <= "1111111111";
                when x"128E" => data <= "1111111111";
                when x"128F" => data <= "1111111111";
                when x"1290" => data <= "1111111111";
                when x"1291" => data <= "1111111111";
                when x"1292" => data <= "1111111111";
                when x"1293" => data <= "1111111111";
                when x"1294" => data <= "1111111111";
                when x"1295" => data <= "1111111111";
                when x"1296" => data <= "1111111111";
                when x"1297" => data <= "1111111111";
                when x"1298" => data <= "1111111111";
                when x"1299" => data <= "1111111111";
                when x"129A" => data <= "1111111111";
                when x"129B" => data <= "1111111111";
                when x"129C" => data <= "1111111111";
                when x"129D" => data <= "1111111111";
                when x"129E" => data <= "1111111111";
                when x"129F" => data <= "1111111111";
                when x"12A0" => data <= "1111111111";
                when x"12A1" => data <= "1111111111";
                when x"12A2" => data <= "1111111111";
                when x"12A3" => data <= "1111111111";
                when x"12A4" => data <= "1111111111";
                when x"12A5" => data <= "1111111111";
                when x"12A6" => data <= "1111111111";
                when x"12A7" => data <= "1111111111";
                when x"12A8" => data <= "1111111111";
                when x"12A9" => data <= "1111111111";
                when x"12AA" => data <= "1111111111";
                when x"12AB" => data <= "1111111111";
                when x"12AC" => data <= "0000100100";
                when x"12AD" => data <= "1111111111";
                when x"12AE" => data <= "1111111111";
                when x"12AF" => data <= "1111111111";
                when x"12B0" => data <= "1111111111";
                when x"12B1" => data <= "1111111111";
                when x"12B2" => data <= "1111111111";
                when x"12B3" => data <= "1111111111";
                when x"12B4" => data <= "1111111111";
                when x"12B5" => data <= "1111111111";
                when x"12B6" => data <= "1111111111";
                when x"12B7" => data <= "1111111111";
                when x"12B8" => data <= "1111111111";
                when x"12B9" => data <= "1111111111";
                when x"12BA" => data <= "1111111111";
                when x"12BB" => data <= "1111111111";
                when x"12BC" => data <= "1111111111";
                when x"12BD" => data <= "1111111111";
                when x"12BE" => data <= "1111111111";
                when x"12BF" => data <= "1111111111";
                when x"12C0" => data <= "1111111111";
                when x"12C1" => data <= "1111111111";
                when x"12C2" => data <= "1111111111";
                when x"12C3" => data <= "1111111111";
                when x"12C4" => data <= "1111111111";
                when x"12C5" => data <= "1111111111";
                when x"12C6" => data <= "1111111111";
                when x"12C7" => data <= "1111111111";
                when x"12C8" => data <= "1111111111";
                when x"12C9" => data <= "1111111111";
                when x"12CA" => data <= "1111111111";
                when x"12CB" => data <= "1111111111";
                when x"12CC" => data <= "1111111111";
                when x"12CD" => data <= "1111111111";
                when x"12CE" => data <= "1111111111";
                when x"12CF" => data <= "1111111111";
                when x"12D0" => data <= "1111111111";
                when x"12D1" => data <= "1111111111";
                when x"12D2" => data <= "1111111111";
                when x"12D3" => data <= "1111111111";
                when x"12D4" => data <= "1111111111";
                when x"12D5" => data <= "1111111111";
                when x"12D6" => data <= "1111111111";
                when x"12D7" => data <= "1111111111";
                when x"12D8" => data <= "1111111111";
                when x"12D9" => data <= "1111111111";
                when x"12DA" => data <= "1111111111";
                when x"12DB" => data <= "1111111111";
                when x"12DC" => data <= "1111111111";
                when x"12DD" => data <= "1111111111";
                when x"12DE" => data <= "1111111111";
                when x"12DF" => data <= "1111111111";
                when x"12E0" => data <= "1111111111";
                when x"12E1" => data <= "1111111111";
                when x"12E2" => data <= "1111111111";
                when x"12E3" => data <= "1111111111";
                when x"12E4" => data <= "1111111111";
                when x"12E5" => data <= "1111111111";
                when x"12E6" => data <= "1111111111";
                when x"12E7" => data <= "1111111111";
                when x"12E8" => data <= "1111111111";
                when x"12E9" => data <= "1011101001";
                when x"12EA" => data <= "1111111111";
                when x"12EB" => data <= "1111111111";
                when x"12EC" => data <= "1111111111";
                when x"12ED" => data <= "1111111111";
                when x"12EE" => data <= "1111111111";
                when x"12EF" => data <= "1111111111";
                when x"12F0" => data <= "1111111111";
                when x"12F1" => data <= "1111111111";
                when x"12F2" => data <= "1111111111";
                when x"12F3" => data <= "1111111111";
                when x"12F4" => data <= "1111111111";
                when x"12F5" => data <= "1111111111";
                when x"12F6" => data <= "1111111111";
                when x"12F7" => data <= "1111111111";
                when x"12F8" => data <= "1111111111";
                when x"12F9" => data <= "1111111111";
                when x"12FA" => data <= "1111111111";
                when x"12FB" => data <= "1111111111";
                when x"12FC" => data <= "1111111111";
                when x"12FD" => data <= "1111111111";
                when x"12FE" => data <= "1111111111";
                when x"12FF" => data <= "1111111111";
                when x"1300" => data <= "1111111111";
                when x"1301" => data <= "1111111111";
                when x"1302" => data <= "1111111111";
                when x"1303" => data <= "1111111111";
                when x"1304" => data <= "1111111111";
                when x"1305" => data <= "1111111111";
                when x"1306" => data <= "1111111111";
                when x"1307" => data <= "1111111111";
                when x"1308" => data <= "1111111111";
                when x"1309" => data <= "1111111111";
                when x"130A" => data <= "1111111111";
                when x"130B" => data <= "1111111111";
                when x"130C" => data <= "1111111111";
                when x"130D" => data <= "1111111111";
                when x"130E" => data <= "1111111111";
                when x"130F" => data <= "1111111111";
                when x"1310" => data <= "1111111111";
                when x"1311" => data <= "1111111111";
                when x"1312" => data <= "1111111111";
                when x"1313" => data <= "1111111111";
                when x"1314" => data <= "1111111111";
                when x"1315" => data <= "1111111111";
                when x"1316" => data <= "1111111111";
                when x"1317" => data <= "1111111111";
                when x"1318" => data <= "1111111111";
                when x"1319" => data <= "1111111111";
                when x"131A" => data <= "1111111111";
                when x"131B" => data <= "1111111111";
                when x"131C" => data <= "1111111111";
                when x"131D" => data <= "1111111111";
                when x"131E" => data <= "1111111111";
                when x"131F" => data <= "1111111111";
                when x"1320" => data <= "1111111111";
                when x"1321" => data <= "1111111111";
                when x"1322" => data <= "1111111111";
                when x"1323" => data <= "1111111111";
                when x"1324" => data <= "1111111111";
                when x"1325" => data <= "1111111111";
                when x"1326" => data <= "1111111111";
                when x"1327" => data <= "1111111111";
                when x"1328" => data <= "1111111111";
                when x"1329" => data <= "1111111111";
                when x"132A" => data <= "1111111111";
                when x"132B" => data <= "1111111111";
                when x"132C" => data <= "1111111111";
                when x"132D" => data <= "1111111111";
                when x"132E" => data <= "1111111111";
                when x"132F" => data <= "1111111111";
                when x"1330" => data <= "1111111111";
                when x"1331" => data <= "1111111111";
                when x"1332" => data <= "1111111111";
                when x"1333" => data <= "1111111111";
                when x"1334" => data <= "1111111111";
                when x"1335" => data <= "1111111111";
                when x"1336" => data <= "1111111111";
                when x"1337" => data <= "1111111111";
                when x"1338" => data <= "1111111111";
                when x"1339" => data <= "1111111111";
                when x"133A" => data <= "1111111111";
                when x"133B" => data <= "1111111111";
                when x"133C" => data <= "1111111111";
                when x"133D" => data <= "1111111111";
                when x"133E" => data <= "1111111111";
                when x"133F" => data <= "1111111111";
                when x"1340" => data <= "1111111111";
                when x"1341" => data <= "1111111111";
                when x"1342" => data <= "1111111111";
                when x"1343" => data <= "1111111111";
                when x"1344" => data <= "1111111111";
                when x"1345" => data <= "1000001000";
                when x"1346" => data <= "1111111111";
                when x"1347" => data <= "1111111111";
                when x"1348" => data <= "1111111111";
                when x"1349" => data <= "1111111111";
                when x"134A" => data <= "1111111111";
                when x"134B" => data <= "1111111111";
                when x"134C" => data <= "1111111111";
                when x"134D" => data <= "1111111111";
                when x"134E" => data <= "1111111111";
                when x"134F" => data <= "1111111111";
                when x"1350" => data <= "1111111111";
                when x"1351" => data <= "1111111111";
                when x"1352" => data <= "1111111111";
                when x"1353" => data <= "1111111111";
                when x"1354" => data <= "1111111111";
                when x"1355" => data <= "1111111111";
                when x"1356" => data <= "1111111111";
                when x"1357" => data <= "1111111111";
                when x"1358" => data <= "1111111111";
                when x"1359" => data <= "1111111111";
                when x"135A" => data <= "1111111111";
                when x"135B" => data <= "1111111111";
                when x"135C" => data <= "1111111111";
                when x"135D" => data <= "1111111111";
                when x"135E" => data <= "1111111111";
                when x"135F" => data <= "1000001000";
                when x"1360" => data <= "1111111111";
                when x"1361" => data <= "1111111111";
                when x"1362" => data <= "1111111111";
                when x"1363" => data <= "1111111111";
                when x"1364" => data <= "1111111111";
                when x"1365" => data <= "1111111111";
                when x"1366" => data <= "1111111111";
                when x"1367" => data <= "1111111111";
                when x"1368" => data <= "1111111111";
                when x"1369" => data <= "1111111111";
                when x"136A" => data <= "1111111111";
                when x"136B" => data <= "1111111111";
                when x"136C" => data <= "1111111111";
                when x"136D" => data <= "1111111111";
                when x"136E" => data <= "1111111111";
                when x"136F" => data <= "1111111111";
                when x"1370" => data <= "1111111111";
                when x"1371" => data <= "1111111111";
                when x"1372" => data <= "1111111111";
                when x"1373" => data <= "1111111111";
                when x"1374" => data <= "1111111111";
                when x"1375" => data <= "1111111111";
                when x"1376" => data <= "1111111111";
                when x"1377" => data <= "1111111111";
                when x"1378" => data <= "1111111111";
                when x"1379" => data <= "1111111111";
                when x"137A" => data <= "1111111111";
                when x"137B" => data <= "1111111111";
                when x"137C" => data <= "1111111111";
                when x"137D" => data <= "0101101101";
                when x"137E" => data <= "1111111111";
                when x"137F" => data <= "1111111111";
                when x"1380" => data <= "1111111111";
                when x"1381" => data <= "1111111111";
                when x"1382" => data <= "1111111111";
                when x"1383" => data <= "1111111111";
                when x"1384" => data <= "1111111111";
                when x"1385" => data <= "1111111111";
                when x"1386" => data <= "1111111111";
                when x"1387" => data <= "1111111111";
                when x"1388" => data <= "1111111111";
                when x"1389" => data <= "1111111111";
                when x"138A" => data <= "1111111111";
                when x"138B" => data <= "1111111111";
                when x"138C" => data <= "1111111111";
                when x"138D" => data <= "1111111111";
                when x"138E" => data <= "1111111111";
                when x"138F" => data <= "1111111111";
                when x"1390" => data <= "1111111111";
                when x"1391" => data <= "1111111111";
                when x"1392" => data <= "1111111111";
                when x"1393" => data <= "1111111111";
                when x"1394" => data <= "1111111111";
                when x"1395" => data <= "1111111111";
                when x"1396" => data <= "1111111111";
                when x"1397" => data <= "1111111111";
                when x"1398" => data <= "1111111111";
                when x"1399" => data <= "1111111111";
                when x"139A" => data <= "1111111111";
                when x"139B" => data <= "1111111111";
                when x"139C" => data <= "1111111111";
                when x"139D" => data <= "1111111111";
                when x"139E" => data <= "1111111111";
                when x"139F" => data <= "1111111111";
                when x"13A0" => data <= "1111111111";
                when x"13A1" => data <= "1111111111";
                when x"13A2" => data <= "1111111111";
                when x"13A3" => data <= "1111111111";
                when x"13A4" => data <= "1111111111";
                when x"13A5" => data <= "1111111111";
                when x"13A6" => data <= "1111111111";
                when x"13A7" => data <= "1111111111";
                when x"13A8" => data <= "1111111111";
                when x"13A9" => data <= "1111111111";
                when x"13AA" => data <= "1111111111";
                when x"13AB" => data <= "1111111111";
                when x"13AC" => data <= "1111111111";
                when x"13AD" => data <= "1111111111";
                when x"13AE" => data <= "1111111111";
                when x"13AF" => data <= "1111111111";
                when x"13B0" => data <= "1111111111";
                when x"13B1" => data <= "1111111111";
                when x"13B2" => data <= "1111111111";
                when x"13B3" => data <= "1111111111";
                when x"13B4" => data <= "1111111111";
                when x"13B5" => data <= "1111111111";
                when x"13B6" => data <= "1111111111";
                when x"13B7" => data <= "1111111111";
                when x"13B8" => data <= "1111111111";
                when x"13B9" => data <= "1111111111";
                when x"13BA" => data <= "1111111111";
                when x"13BB" => data <= "1111111111";
                when x"13BC" => data <= "1111111111";
                when x"13BD" => data <= "1111111111";
                when x"13BE" => data <= "1111111111";
                when x"13BF" => data <= "1111111111";
                when x"13C0" => data <= "1111111111";
                when x"13C1" => data <= "1111111111";
                when x"13C2" => data <= "1111111111";
                when x"13C3" => data <= "1111111111";
                when x"13C4" => data <= "1111111111";
                when x"13C5" => data <= "1111111111";
                when x"13C6" => data <= "1111111111";
                when x"13C7" => data <= "1111111111";
                when x"13C8" => data <= "1111111111";
                when x"13C9" => data <= "1111111111";
                when x"13CA" => data <= "1111111111";
                when x"13CB" => data <= "1111111111";
                when x"13CC" => data <= "1111111111";
                when x"13CD" => data <= "1111111111";
                when x"13CE" => data <= "1111111111";
                when x"13CF" => data <= "1111111111";
                when x"13D0" => data <= "1000001000";
                when x"13D1" => data <= "1111111111";
                when x"13D2" => data <= "1111111111";
                when x"13D3" => data <= "0001111011";
                when x"13D4" => data <= "1111111111";
                when x"13D5" => data <= "1111111111";
                when x"13D6" => data <= "1111111111";
                when x"13D7" => data <= "1111111111";
                when x"13D8" => data <= "1111111111";
                when x"13D9" => data <= "1111111111";
                when x"13DA" => data <= "1111111111";
                when x"13DB" => data <= "1111111111";
                when x"13DC" => data <= "1111111111";
                when x"13DD" => data <= "1000001000";
                when x"13DE" => data <= "1111111111";
                when x"13DF" => data <= "1111111111";
                when x"13E0" => data <= "1111111111";
                when x"13E1" => data <= "1111111111";
                when x"13E2" => data <= "1111111111";
                when x"13E3" => data <= "1111111111";
                when x"13E4" => data <= "1111111111";
                when x"13E5" => data <= "1111111111";
                when x"13E6" => data <= "1111111111";
                when x"13E7" => data <= "1111111111";
                when x"13E8" => data <= "1000001000";
                when x"13E9" => data <= "1111111111";
                when x"13EA" => data <= "1111111111";
                when x"13EB" => data <= "1111111111";
                when x"13EC" => data <= "1111111111";
                when x"13ED" => data <= "1111111111";
                when x"13EE" => data <= "1111111111";
                when x"13EF" => data <= "1111111111";
                when x"13F0" => data <= "1111111111";
                when x"13F1" => data <= "1111111111";
                when x"13F2" => data <= "1111111111";
                when x"13F3" => data <= "1111111111";
                when x"13F4" => data <= "1111111111";
                when x"13F5" => data <= "1111111111";
                when x"13F6" => data <= "1111111111";
                when x"13F7" => data <= "1111111111";
                when x"13F8" => data <= "1111111111";
                when x"13F9" => data <= "1111111111";
                when x"13FA" => data <= "1111111111";
                when x"13FB" => data <= "1111111111";
                when x"13FC" => data <= "1111111111";
                when x"13FD" => data <= "1111111111";
                when x"13FE" => data <= "1111111111";
                when x"13FF" => data <= "1111111111";
                when x"1400" => data <= "1111111111";
                when x"1401" => data <= "1111111111";
                when x"1402" => data <= "1111111111";
                when x"1403" => data <= "1111111111";
                when x"1404" => data <= "1111111111";
                when x"1405" => data <= "1111111111";
                when x"1406" => data <= "1111111111";
                when x"1407" => data <= "1111111111";
                when x"1408" => data <= "1111111111";
                when x"1409" => data <= "1111111111";
                when x"140A" => data <= "1111111111";
                when x"140B" => data <= "1111111111";
                when x"140C" => data <= "1111111111";
                when x"140D" => data <= "1111111111";
                when x"140E" => data <= "1111111111";
                when x"140F" => data <= "1111111111";
                when x"1410" => data <= "1111111111";
                when x"1411" => data <= "1111111111";
                when x"1412" => data <= "1111111111";
                when x"1413" => data <= "1111111111";
                when x"1414" => data <= "1111111111";
                when x"1415" => data <= "1111111111";
                when x"1416" => data <= "1111111111";
                when x"1417" => data <= "1111111111";
                when x"1418" => data <= "1111111111";
                when x"1419" => data <= "1111111111";
                when x"141A" => data <= "1111111111";
                when x"141B" => data <= "1111111111";
                when x"141C" => data <= "1111111111";
                when x"141D" => data <= "1111111111";
                when x"141E" => data <= "1111111111";
                when x"141F" => data <= "1111111111";
                when x"1420" => data <= "1111111111";
                when x"1421" => data <= "1111111111";
                when x"1422" => data <= "1111111111";
                when x"1423" => data <= "1111111111";
                when x"1424" => data <= "1111111111";
                when x"1425" => data <= "1111111111";
                when x"1426" => data <= "1111111111";
                when x"1427" => data <= "1111111111";
                when x"1428" => data <= "1111111111";
                when x"1429" => data <= "1111111111";
                when x"142A" => data <= "1111111111";
                when x"142B" => data <= "1111111111";
                when x"142C" => data <= "1111111111";
                when x"142D" => data <= "1111111111";
                when x"142E" => data <= "1111111111";
                when x"142F" => data <= "1111111111";
                when x"1430" => data <= "1111111111";
                when x"1431" => data <= "1111111111";
                when x"1432" => data <= "1111111111";
                when x"1433" => data <= "1111111111";
                when x"1434" => data <= "1111111111";
                when x"1435" => data <= "1111111111";
                when x"1436" => data <= "1111111111";
                when x"1437" => data <= "1111111111";
                when x"1438" => data <= "1111111111";
                when x"1439" => data <= "1111111111";
                when x"143A" => data <= "1111111111";
                when x"143B" => data <= "1111111111";
                when x"143C" => data <= "1111111111";
                when x"143D" => data <= "1111111111";
                when x"143E" => data <= "1111111111";
                when x"143F" => data <= "1111111111";
                when x"1440" => data <= "1111111111";
                when x"1441" => data <= "1111111111";
                when x"1442" => data <= "1111111111";
                when x"1443" => data <= "1111111111";
                when x"1444" => data <= "1111111111";
                when x"1445" => data <= "1111111111";
                when x"1446" => data <= "1111111111";
                when x"1447" => data <= "1111111111";
                when x"1448" => data <= "1111111111";
                when x"1449" => data <= "1111111111";
                when x"144A" => data <= "1111111111";
                when x"144B" => data <= "1111111111";
                when x"144C" => data <= "1111111111";
                when x"144D" => data <= "1111111111";
                when x"144E" => data <= "1111111111";
                when x"144F" => data <= "1111111111";
                when x"1450" => data <= "1111111111";
                when x"1451" => data <= "1111111111";
                when x"1452" => data <= "1111111111";
                when x"1453" => data <= "1111111111";
                when x"1454" => data <= "1111111111";
                when x"1455" => data <= "1111111111";
                when x"1456" => data <= "1111111111";
                when x"1457" => data <= "1111111111";
                when x"1458" => data <= "1111111111";
                when x"1459" => data <= "1111111111";
                when x"145A" => data <= "1111111111";
                when x"145B" => data <= "1111111111";
                when x"145C" => data <= "1111111111";
                when x"145D" => data <= "1111111111";
                when x"145E" => data <= "1111111111";
                when x"145F" => data <= "1111111111";
                when x"1460" => data <= "1111111111";
                when x"1461" => data <= "1111111111";
                when x"1462" => data <= "1111111111";
                when x"1463" => data <= "1111111111";
                when x"1464" => data <= "1111111111";
                when x"1465" => data <= "1111111111";
                when x"1466" => data <= "1111111111";
                when x"1467" => data <= "1111111111";
                when x"1468" => data <= "1111111111";
                when x"1469" => data <= "0101101101";
                when x"146A" => data <= "1111111111";
                when x"146B" => data <= "1111111111";
                when x"146C" => data <= "1111111111";
                when x"146D" => data <= "1111111111";
                when x"146E" => data <= "1111111111";
                when x"146F" => data <= "1111111111";
                when x"1470" => data <= "1111111111";
                when x"1471" => data <= "1111111111";
                when x"1472" => data <= "1111111111";
                when x"1473" => data <= "1111111111";
                when x"1474" => data <= "1111111111";
                when x"1475" => data <= "1111111111";
                when x"1476" => data <= "1111111111";
                when x"1477" => data <= "1111111111";
                when x"1478" => data <= "1111111111";
                when x"1479" => data <= "1111111111";
                when x"147A" => data <= "1111111111";
                when x"147B" => data <= "1111111111";
                when x"147C" => data <= "1111111111";
                when x"147D" => data <= "1111111111";
                when x"147E" => data <= "1111111111";
                when x"147F" => data <= "1111111111";
                when x"1480" => data <= "1111111111";
                when x"1481" => data <= "1111111111";
                when x"1482" => data <= "1111111111";
                when x"1483" => data <= "1111111111";
                when x"1484" => data <= "1111111111";
                when x"1485" => data <= "1111111111";
                when x"1486" => data <= "1111111111";
                when x"1487" => data <= "1111111111";
                when x"1488" => data <= "1111111111";
                when x"1489" => data <= "1111111111";
                when x"148A" => data <= "1111111111";
                when x"148B" => data <= "1111111111";
                when x"148C" => data <= "1111111111";
                when x"148D" => data <= "1111111111";
                when x"148E" => data <= "1111111111";
                when x"148F" => data <= "1111111111";
                when x"1490" => data <= "1111111111";
                when x"1491" => data <= "1111111111";
                when x"1492" => data <= "1111111111";
                when x"1493" => data <= "1111111111";
                when x"1494" => data <= "1111111111";
                when x"1495" => data <= "1111111111";
                when x"1496" => data <= "1111111111";
                when x"1497" => data <= "1111111111";
                when x"1498" => data <= "1111111111";
                when x"1499" => data <= "1111111111";
                when x"149A" => data <= "1111111111";
                when x"149B" => data <= "1111111111";
                when x"149C" => data <= "1111111111";
                when x"149D" => data <= "1111111111";
                when x"149E" => data <= "1111111111";
                when x"149F" => data <= "1111111111";
                when x"14A0" => data <= "1111111111";
                when x"14A1" => data <= "1111111111";
                when x"14A2" => data <= "1111111111";
                when x"14A3" => data <= "1111111111";
                when x"14A4" => data <= "1111111111";
                when x"14A5" => data <= "1111111111";
                when x"14A6" => data <= "1111111111";
                when x"14A7" => data <= "1111111111";
                when x"14A8" => data <= "1111111111";
                when x"14A9" => data <= "1111111111";
                when x"14AA" => data <= "1111111111";
                when x"14AB" => data <= "1111111111";
                when x"14AC" => data <= "1111111111";
                when x"14AD" => data <= "1111111111";
                when x"14AE" => data <= "1111111111";
                when x"14AF" => data <= "1111111111";
                when x"14B0" => data <= "1111111111";
                when x"14B1" => data <= "1111111111";
                when x"14B2" => data <= "1111111111";
                when x"14B3" => data <= "1111111111";
                when x"14B4" => data <= "1111111111";
                when x"14B5" => data <= "1111111111";
                when x"14B6" => data <= "1111111111";
                when x"14B7" => data <= "1111111111";
                when x"14B8" => data <= "1111111111";
                when x"14B9" => data <= "1111111111";
                when x"14BA" => data <= "1111111111";
                when x"14BB" => data <= "1111111111";
                when x"14BC" => data <= "1111111111";
                when x"14BD" => data <= "1111111111";
                when x"14BE" => data <= "1111111111";
                when x"14BF" => data <= "1111111111";
                when x"14C0" => data <= "1111111111";
                when x"14C1" => data <= "1111111111";
                when x"14C2" => data <= "1111111111";
                when x"14C3" => data <= "1111111111";
                when x"14C4" => data <= "1111111111";
                when x"14C5" => data <= "1111111111";
                when x"14C6" => data <= "1111111111";
                when x"14C7" => data <= "1111111111";
                when x"14C8" => data <= "1111111111";
                when x"14C9" => data <= "1111111111";
                when x"14CA" => data <= "1111111111";
                when x"14CB" => data <= "1111111111";
                when x"14CC" => data <= "1111111111";
                when x"14CD" => data <= "1111111111";
                when x"14CE" => data <= "1111111111";
                when x"14CF" => data <= "1111111111";
                when x"14D0" => data <= "1111111111";
                when x"14D1" => data <= "1111111111";
                when x"14D2" => data <= "1111111111";
                when x"14D3" => data <= "1111111111";
                when x"14D4" => data <= "1111111111";
                when x"14D5" => data <= "1111111111";
                when x"14D6" => data <= "1111111111";
                when x"14D7" => data <= "1111111111";
                when x"14D8" => data <= "1111111111";
                when x"14D9" => data <= "1111111111";
                when x"14DA" => data <= "1111111111";
                when x"14DB" => data <= "1111111111";
                when x"14DC" => data <= "1111111111";
                when x"14DD" => data <= "1111111111";
                when x"14DE" => data <= "1111111111";
                when x"14DF" => data <= "1111111111";
                when x"14E0" => data <= "1111111111";
                when x"14E1" => data <= "1111111111";
                when x"14E2" => data <= "1111111111";
                when x"14E3" => data <= "1111111111";
                when x"14E4" => data <= "1111111111";
                when x"14E5" => data <= "1111111111";
                when x"14E6" => data <= "1111111111";
                when x"14E7" => data <= "1111111111";
                when x"14E8" => data <= "1111111111";
                when x"14E9" => data <= "1111111111";
                when x"14EA" => data <= "1111111111";
                when x"14EB" => data <= "1111111111";
                when x"14EC" => data <= "1111111111";
                when x"14ED" => data <= "1111111111";
                when x"14EE" => data <= "1111111111";
                when x"14EF" => data <= "1111111111";
                when x"14F0" => data <= "1111111111";
                when x"14F1" => data <= "1111111111";
                when x"14F2" => data <= "1111111111";
                when x"14F3" => data <= "1111111111";
                when x"14F4" => data <= "1111111111";
                when x"14F5" => data <= "1111111111";
                when x"14F6" => data <= "1111111111";
                when x"14F7" => data <= "1111111111";
                when x"14F8" => data <= "1111111111";
                when x"14F9" => data <= "1111111111";
                when x"14FA" => data <= "1111111111";
                when x"14FB" => data <= "1111111111";
                when x"14FC" => data <= "1111111111";
                when x"14FD" => data <= "1111111111";
                when x"14FE" => data <= "1111111111";
                when x"14FF" => data <= "1111111111";
                when x"1500" => data <= "1111111111";
                when x"1501" => data <= "1111111111";
                when x"1502" => data <= "1111111111";
                when x"1503" => data <= "1111111111";
                when x"1504" => data <= "1111111111";
                when x"1505" => data <= "1111111111";
                when x"1506" => data <= "1111111111";
                when x"1507" => data <= "1111111111";
                when x"1508" => data <= "1111111111";
                when x"1509" => data <= "1111111111";
                when x"150A" => data <= "1111111111";
                when x"150B" => data <= "1111111111";
                when x"150C" => data <= "1111111111";
                when x"150D" => data <= "1111111111";
                when x"150E" => data <= "1111111111";
                when x"150F" => data <= "1111111111";
                when x"1510" => data <= "1111111111";
                when x"1511" => data <= "1111111111";
                when x"1512" => data <= "1111111111";
                when x"1513" => data <= "1111111111";
                when x"1514" => data <= "1111111111";
                when x"1515" => data <= "1111111111";
                when x"1516" => data <= "1111111111";
                when x"1517" => data <= "1111111111";
                when x"1518" => data <= "1111111111";
                when x"1519" => data <= "1111111111";
                when x"151A" => data <= "1111111111";
                when x"151B" => data <= "1111111111";
                when x"151C" => data <= "1111111111";
                when x"151D" => data <= "1111111111";
                when x"151E" => data <= "1111111111";
                when x"151F" => data <= "1111111111";
                when x"1520" => data <= "1111111111";
                when x"1521" => data <= "1111111111";
                when x"1522" => data <= "1111111111";
                when x"1523" => data <= "1111111111";
                when x"1524" => data <= "0101011000";
                when x"1525" => data <= "1111111111";
                when x"1526" => data <= "1111111111";
                when x"1527" => data <= "1111111111";
                when x"1528" => data <= "1111111111";
                when x"1529" => data <= "1111111111";
                when x"152A" => data <= "1111111111";
                when x"152B" => data <= "1111111111";
                when x"152C" => data <= "1111111111";
                when x"152D" => data <= "1111111111";
                when x"152E" => data <= "1111111111";
                when x"152F" => data <= "1111111111";
                when x"1530" => data <= "1111111111";
                when x"1531" => data <= "1111111111";
                when x"1532" => data <= "1111111111";
                when x"1533" => data <= "1111111111";
                when x"1534" => data <= "1111111111";
                when x"1535" => data <= "1111111111";
                when x"1536" => data <= "1111111111";
                when x"1537" => data <= "1111111111";
                when x"1538" => data <= "1111111111";
                when x"1539" => data <= "1111111111";
                when x"153A" => data <= "1111111111";
                when x"153B" => data <= "1111111111";
                when x"153C" => data <= "1111111111";
                when x"153D" => data <= "1111111111";
                when x"153E" => data <= "1111111111";
                when x"153F" => data <= "1111111111";
                when x"1540" => data <= "1111111111";
                when x"1541" => data <= "1111111111";
                when x"1542" => data <= "1111111111";
                when x"1543" => data <= "1111111111";
                when x"1544" => data <= "1111111111";
                when x"1545" => data <= "1111111111";
                when x"1546" => data <= "1111111111";
                when x"1547" => data <= "1111111111";
                when x"1548" => data <= "1111111111";
                when x"1549" => data <= "1111111111";
                when x"154A" => data <= "1111111111";
                when x"154B" => data <= "1111111111";
                when x"154C" => data <= "1111111111";
                when x"154D" => data <= "1111111111";
                when x"154E" => data <= "1111111111";
                when x"154F" => data <= "1111111111";
                when x"1550" => data <= "1111111111";
                when x"1551" => data <= "1111111111";
                when x"1552" => data <= "1111111111";
                when x"1553" => data <= "1111111111";
                when x"1554" => data <= "1111111111";
                when x"1555" => data <= "1111111111";
                when x"1556" => data <= "1111111111";
                when x"1557" => data <= "1111111111";
                when x"1558" => data <= "1111111111";
                when x"1559" => data <= "1111111111";
                when x"155A" => data <= "1111111111";
                when x"155B" => data <= "1111111111";
                when x"155C" => data <= "1111111111";
                when x"155D" => data <= "1111111111";
                when x"155E" => data <= "1000111101";
                when x"155F" => data <= "1111111111";
                when x"1560" => data <= "1111111111";
                when x"1561" => data <= "1111111111";
                when x"1562" => data <= "1111111111";
                when x"1563" => data <= "1111111111";
                when x"1564" => data <= "1111111111";
                when x"1565" => data <= "1111111111";
                when x"1566" => data <= "1111111111";
                when x"1567" => data <= "1111111111";
                when x"1568" => data <= "1111111111";
                when x"1569" => data <= "1111111111";
                when x"156A" => data <= "1111111111";
                when x"156B" => data <= "1111111111";
                when x"156C" => data <= "1111111111";
                when x"156D" => data <= "1111111111";
                when x"156E" => data <= "1111111111";
                when x"156F" => data <= "1111111111";
                when x"1570" => data <= "1111111111";
                when x"1571" => data <= "1111111111";
                when x"1572" => data <= "1111111111";
                when x"1573" => data <= "1111111111";
                when x"1574" => data <= "1111111111";
                when x"1575" => data <= "1111111111";
                when x"1576" => data <= "1111111111";
                when x"1577" => data <= "1111111111";
                when x"1578" => data <= "1111111111";
                when x"1579" => data <= "1111111111";
                when x"157A" => data <= "1111111111";
                when x"157B" => data <= "1111111111";
                when x"157C" => data <= "1111111111";
                when x"157D" => data <= "1111111111";
                when x"157E" => data <= "1111111111";
                when x"157F" => data <= "1111111111";
                when x"1580" => data <= "1111111111";
                when x"1581" => data <= "1111111111";
                when x"1582" => data <= "1111111111";
                when x"1583" => data <= "1111111111";
                when x"1584" => data <= "1111111111";
                when x"1585" => data <= "1111111111";
                when x"1586" => data <= "1111111111";
                when x"1587" => data <= "1111111111";
                when x"1588" => data <= "1111111111";
                when x"1589" => data <= "1111111111";
                when x"158A" => data <= "1111111111";
                when x"158B" => data <= "1111111111";
                when x"158C" => data <= "1111111111";
                when x"158D" => data <= "1111111111";
                when x"158E" => data <= "1111111111";
                when x"158F" => data <= "1111111111";
                when x"1590" => data <= "1111111111";
                when x"1591" => data <= "1111111111";
                when x"1592" => data <= "1111111111";
                when x"1593" => data <= "1111111111";
                when x"1594" => data <= "1111111111";
                when x"1595" => data <= "1111111111";
                when x"1596" => data <= "1111111111";
                when x"1597" => data <= "1111111111";
                when x"1598" => data <= "1111111111";
                when x"1599" => data <= "1111111111";
                when x"159A" => data <= "1111111111";
                when x"159B" => data <= "1111111111";
                when x"159C" => data <= "1111111111";
                when x"159D" => data <= "1111111111";
                when x"159E" => data <= "1111111111";
                when x"159F" => data <= "1111111111";
                when x"15A0" => data <= "1111111111";
                when x"15A1" => data <= "1111111111";
                when x"15A2" => data <= "1111111111";
                when x"15A3" => data <= "1111111111";
                when x"15A4" => data <= "1111111111";
                when x"15A5" => data <= "1111111111";
                when x"15A6" => data <= "1111111111";
                when x"15A7" => data <= "1111111111";
                when x"15A8" => data <= "1111111111";
                when x"15A9" => data <= "1111111111";
                when x"15AA" => data <= "1111111111";
                when x"15AB" => data <= "1111111111";
                when x"15AC" => data <= "1111111111";
                when x"15AD" => data <= "1111111111";
                when x"15AE" => data <= "1111111111";
                when x"15AF" => data <= "1111111111";
                when x"15B0" => data <= "1111111111";
                when x"15B1" => data <= "1111111111";
                when x"15B2" => data <= "1111111111";
                when x"15B3" => data <= "1111111111";
                when x"15B4" => data <= "1111111111";
                when x"15B5" => data <= "1111111111";
                when x"15B6" => data <= "1111111111";
                when x"15B7" => data <= "1111111111";
                when x"15B8" => data <= "1111111111";
                when x"15B9" => data <= "1111111111";
                when x"15BA" => data <= "1111111111";
                when x"15BB" => data <= "1111111111";
                when x"15BC" => data <= "1111111111";
                when x"15BD" => data <= "1111111111";
                when x"15BE" => data <= "1111111111";
                when x"15BF" => data <= "1111111111";
                when x"15C0" => data <= "1111111111";
                when x"15C1" => data <= "1111111111";
                when x"15C2" => data <= "1111111111";
                when x"15C3" => data <= "1111111111";
                when x"15C4" => data <= "1111111111";
                when x"15C5" => data <= "1111111111";
                when x"15C6" => data <= "1111111111";
                when x"15C7" => data <= "1111111111";
                when x"15C8" => data <= "1111111111";
                when x"15C9" => data <= "1111111111";
                when x"15CA" => data <= "1111111111";
                when x"15CB" => data <= "1111111111";
                when x"15CC" => data <= "1111111111";
                when x"15CD" => data <= "1111111111";
                when x"15CE" => data <= "1111111111";
                when x"15CF" => data <= "1111111111";
                when x"15D0" => data <= "1111111111";
                when x"15D1" => data <= "1111111111";
                when x"15D2" => data <= "1111111111";
                when x"15D3" => data <= "1111111111";
                when x"15D4" => data <= "1111111111";
                when x"15D5" => data <= "1111111111";
                when x"15D6" => data <= "1111111111";
                when x"15D7" => data <= "1111111111";
                when x"15D8" => data <= "1111111111";
                when x"15D9" => data <= "1111111111";
                when x"15DA" => data <= "1111111111";
                when x"15DB" => data <= "1111111111";
                when x"15DC" => data <= "1111111111";
                when x"15DD" => data <= "1111111111";
                when x"15DE" => data <= "1111111111";
                when x"15DF" => data <= "1111111111";
                when x"15E0" => data <= "1111111111";
                when x"15E1" => data <= "1111111111";
                when x"15E2" => data <= "1111111111";
                when x"15E3" => data <= "1111111111";
                when x"15E4" => data <= "1111111111";
                when x"15E5" => data <= "1111111111";
                when x"15E6" => data <= "1111111111";
                when x"15E7" => data <= "1111111111";
                when x"15E8" => data <= "1111111111";
                when x"15E9" => data <= "1111111111";
                when x"15EA" => data <= "1111111111";
                when x"15EB" => data <= "1111111111";
                when x"15EC" => data <= "1111111111";
                when x"15ED" => data <= "1111111111";
                when x"15EE" => data <= "1111111111";
                when x"15EF" => data <= "1111111111";
                when x"15F0" => data <= "1111111111";
                when x"15F1" => data <= "1111111111";
                when x"15F2" => data <= "1111111111";
                when x"15F3" => data <= "1111111111";
                when x"15F4" => data <= "1111111111";
                when x"15F5" => data <= "1111111111";
                when x"15F6" => data <= "1111111111";
                when x"15F7" => data <= "1111111111";
                when x"15F8" => data <= "1111111111";
                when x"15F9" => data <= "1111111111";
                when x"15FA" => data <= "1111111111";
                when x"15FB" => data <= "1111111111";
                when x"15FC" => data <= "1111111111";
                when x"15FD" => data <= "1111111111";
                when x"15FE" => data <= "1111111111";
                when x"15FF" => data <= "0100000111";
                when x"1600" => data <= "1111111111";
                when x"1601" => data <= "1111111111";
                when x"1602" => data <= "1111111111";
                when x"1603" => data <= "1111111111";
                when x"1604" => data <= "1111111111";
                when x"1605" => data <= "1111111111";
                when x"1606" => data <= "1111111111";
                when x"1607" => data <= "1111111111";
                when x"1608" => data <= "1111111111";
                when x"1609" => data <= "1111111111";
                when x"160A" => data <= "1111111111";
                when x"160B" => data <= "1111111111";
                when x"160C" => data <= "1111111111";
                when x"160D" => data <= "1111111111";
                when x"160E" => data <= "1111111111";
                when x"160F" => data <= "1111111111";
                when x"1610" => data <= "1111111111";
                when x"1611" => data <= "1111111111";
                when x"1612" => data <= "1111111111";
                when x"1613" => data <= "1111111111";
                when x"1614" => data <= "1111111111";
                when x"1615" => data <= "1111111111";
                when x"1616" => data <= "1111111111";
                when x"1617" => data <= "1111111111";
                when x"1618" => data <= "1111111111";
                when x"1619" => data <= "1111111111";
                when x"161A" => data <= "1111111111";
                when x"161B" => data <= "1111111111";
                when x"161C" => data <= "1111111111";
                when x"161D" => data <= "1111111111";
                when x"161E" => data <= "1111111111";
                when x"161F" => data <= "1111111111";
                when x"1620" => data <= "1111111111";
                when x"1621" => data <= "1111111111";
                when x"1622" => data <= "1111111111";
                when x"1623" => data <= "1111111111";
                when x"1624" => data <= "1111111111";
                when x"1625" => data <= "1111111111";
                when x"1626" => data <= "1111111111";
                when x"1627" => data <= "1111111111";
                when x"1628" => data <= "1111111111";
                when x"1629" => data <= "1111111111";
                when x"162A" => data <= "1111111111";
                when x"162B" => data <= "1111111111";
                when x"162C" => data <= "1111111111";
                when x"162D" => data <= "1111111111";
                when x"162E" => data <= "1111111111";
                when x"162F" => data <= "1111111111";
                when x"1630" => data <= "1111111111";
                when x"1631" => data <= "1111111111";
                when x"1632" => data <= "1111111111";
                when x"1633" => data <= "1111111111";
                when x"1634" => data <= "1111111111";
                when x"1635" => data <= "1111111111";
                when x"1636" => data <= "1111111111";
                when x"1637" => data <= "0100010000";
                when x"1638" => data <= "1110000010";
                when x"1639" => data <= "1001000000";
                when x"163A" => data <= "0011010010";
                when x"163B" => data <= "1101010110";
                when x"163C" => data <= "1001000000";
                when x"163D" => data <= "0110101110";
                when x"163E" => data <= "1001000000";
                when x"163F" => data <= "1111011101";
                when x"1640" => data <= "1001000000";
                when x"1641" => data <= "0100100101";
                when x"1642" => data <= "1001000000";
                when x"1643" => data <= "0100100101";
                when x"1644" => data <= "0100100101";
                when x"1645" => data <= "0100100101";
                when x"1646" => data <= "0000000110";
                when x"1647" => data <= "1101010110";
                when x"1648" => data <= "1110110111";
                when x"1649" => data <= "0100100101";
                when x"164A" => data <= "0100100101";
                when x"164B" => data <= "0100010000";
                when x"164C" => data <= "1101010110";
                when x"164D" => data <= "1111101000";
                when x"164E" => data <= "1111011101";
                when x"164F" => data <= "0100100101";
                when x"1650" => data <= "1001000000";
                when x"1651" => data <= "1001000000";
                when x"1652" => data <= "1001110101";
                when x"1653" => data <= "1000011111";
                when x"1654" => data <= "0100100101";
                when x"1655" => data <= "1001000000";
                when x"1656" => data <= "1001000000";
                when x"1657" => data <= "1010100001";
                when x"1658" => data <= "1001000000";
                when x"1659" => data <= "0111000100";
                when x"165A" => data <= "1001000000";
                when x"165B" => data <= "1110000010";
                when x"165C" => data <= "1001000000";
                when x"165D" => data <= "1001110101";
                when x"165E" => data <= "1001000000";
                when x"165F" => data <= "1001000000";
                when x"1660" => data <= "1101010110";
                when x"1661" => data <= "0100100101";
                when x"1662" => data <= "1000101010";
                when x"1663" => data <= "1001000000";
                when x"1664" => data <= "1001000000";
                when x"1665" => data <= "0100100101";
                when x"1666" => data <= "0100010000";
                when x"1667" => data <= "1001000000";
                when x"1668" => data <= "0100100101";
                when x"1669" => data <= "1101010110";
                when x"166A" => data <= "0100010000";
                when x"166B" => data <= "0100010000";
                when x"166C" => data <= "1001000000";
                when x"166D" => data <= "1001000000";
                when x"166E" => data <= "1000101010";
                when x"166F" => data <= "0100100101";
                when x"1670" => data <= "1000000101";
                when x"1671" => data <= "1110011000";
                when x"1672" => data <= "1100010011";
                when x"1673" => data <= "0111101011";
                when x"1674" => data <= "1110011000";
                when x"1675" => data <= "1110011000";
                when x"1676" => data <= "0100111111";
                when x"1677" => data <= "1110101101";
                when x"1678" => data <= "1111110010";
                when x"1679" => data <= "1010001110";
                when x"167A" => data <= "1111110010";
                when x"167B" => data <= "1010111011";
                when x"167C" => data <= "0100001010";
                when x"167D" => data <= "1000110000";
                when x"167E" => data <= "0100111111";
                when x"167F" => data <= "1101111001";
                when x"1680" => data <= "0000101001";
                when x"1681" => data <= "0000101001";
                when x"1682" => data <= "0101010101";
                when x"1683" => data <= "1000000101";
                when x"1684" => data <= "1110101101";
                when x"1685" => data <= "0100111111";
                when x"1686" => data <= "0100001010";
                when x"1687" => data <= "1111000111";
                when x"1688" => data <= "0110000001";
                when x"1689" => data <= "0100111111";
                when x"168A" => data <= "1001011010";
                when x"168B" => data <= "1010111011";
                when x"168C" => data <= "0111011110";
                when x"168D" => data <= "1001011010";
                when x"168E" => data <= "0101010101";
                when x"168F" => data <= "1111110010";
                when x"1690" => data <= "0001000011";
                when x"1691" => data <= "1001101111";
                when x"1692" => data <= "0111011110";
                when x"1693" => data <= "0101010101";
                when x"1694" => data <= "1000000101";
                when x"1695" => data <= "1011100100";
                when x"1696" => data <= "0011001000";
                when x"1697" => data <= "1000000101";
                when x"1698" => data <= "0001110110";
                when x"1699" => data <= "1110101101";
                when x"169A" => data <= "0111011110";
                when x"169B" => data <= "0000101001";
                when x"169C" => data <= "0111101011";
                when x"169D" => data <= "1001100100";
                when x"169E" => data <= "1011011010";
                when x"169F" => data <= "1100011000";
                when x"16A0" => data <= "1011011010";
                when x"16A1" => data <= "0110001010";
                when x"16A2" => data <= "1011101111";
                when x"16A3" => data <= "0110001010";
                when x"16A4" => data <= "0010101001";
                when x"16A5" => data <= "1000111011";
                when x"16A6" => data <= "1011011010";
                when x"16A7" => data <= "0001001000";
                when x"16A8" => data <= "1111001100";
                when x"16A9" => data <= "0111100000";
                when x"16AA" => data <= "0010101001";
                when x"16AB" => data <= "0000100010";
                when x"16AC" => data <= "0110111111";
                when x"16AD" => data <= "1011011010";
                when x"16AE" => data <= "1111111001";
                when x"16AF" => data <= "1011011010";
                when x"16B0" => data <= "0001111101";
                when x"16B1" => data <= "0110001010";
                when x"16B2" => data <= "0000100010";
                when x"16B3" => data <= "0110001010";
                when x"16B4" => data <= "0110111111";
                when x"16B5" => data <= "0110111111";
                when x"16B6" => data <= "0110111111";
                when x"16B7" => data <= "1011101111";
                when x"16B8" => data <= "0110111111";
                when x"16B9" => data <= "1011011010";
                when x"16BA" => data <= "0110111111";
                when x"16BB" => data <= "0110111111";
                when x"16BC" => data <= "0010101001";
                when x"16BD" => data <= "0000100010";
                when x"16BE" => data <= "0110001010";
                when x"16BF" => data <= "0110111111";
                when x"16C0" => data <= "0000010111";
                when x"16C1" => data <= "0110111111";
                when x"16C2" => data <= "1011011010";
                when x"16C3" => data <= "0111010101";
                when x"16C4" => data <= "1011011010";
                when x"16C5" => data <= "1011101111";
                when x"16C6" => data <= "0101011110";
                when x"16C7" => data <= "0110111111";
                when x"16C8" => data <= "0100000001";
                when x"16C9" => data <= "0110111111";
                when x"16CA" => data <= "0111010101";
                when x"16CB" => data <= "1011011010";
                when x"16CC" => data <= "0100000001";
                when x"16CD" => data <= "1010000101";
                when x"16CE" => data <= "0001001000";
                when x"16CF" => data <= "0001001000";
                when x"16D0" => data <= "0110111111";
                when x"16D1" => data <= "0110001010";
                when x"16D2" => data <= "0110001010";
                when x"16D3" => data <= "1101110010";
                when x"16D4" => data <= "0000100010";
                when x"16D5" => data <= "0110111111";
                when x"16D6" => data <= "0010101001";
                when x"16D7" => data <= "0000100010";
                when x"16D8" => data <= "1011011010";
                when x"16D9" => data <= "0110111111";
                when x"16DA" => data <= "0001100111";
                when x"16DB" => data <= "0101000100";
                when x"16DC" => data <= "1011000000";
                when x"16DD" => data <= "1111010110";
                when x"16DE" => data <= "1011110101";
                when x"16DF" => data <= "1100110111";
                when x"16E0" => data <= "0000001101";
                when x"16E1" => data <= "1010101010";
                when x"16E2" => data <= "1000010100";
                when x"16E3" => data <= "1011000000";
                when x"16E4" => data <= "0001100111";
                when x"16E5" => data <= "0110100101";
                when x"16E6" => data <= "0111111010";
                when x"16E7" => data <= "0101000100";
                when x"16E8" => data <= "1011000000";
                when x"16E9" => data <= "1000010100";
                when x"16EA" => data <= "1111010110";
                when x"16EB" => data <= "1011110101";
                when x"16EC" => data <= "0001010010";
                when x"16ED" => data <= "0010110011";
                when x"16EE" => data <= "0000001101";
                when x"16EF" => data <= "0001010010";
                when x"16F0" => data <= "1000100001";
                when x"16F1" => data <= "1111010110";
                when x"16F2" => data <= "0101000100";
                when x"16F3" => data <= "0101000100";
                when x"16F4" => data <= "0101000100";
                when x"16F5" => data <= "0001010010";
                when x"16F6" => data <= "1000100001";
                when x"16F7" => data <= "1011000000";
                when x"16F8" => data <= "0101110001";
                when x"16F9" => data <= "0001010010";
                when x"16FA" => data <= "1111010110";
                when x"16FB" => data <= "0000001101";
                when x"16FC" => data <= "1100110111";
                when x"16FD" => data <= "1011000000";
                when x"16FE" => data <= "1010101010";
                when x"16FF" => data <= "0001100111";
                when x"1700" => data <= "1010011111";
                when x"1701" => data <= "0101000100";
                when x"1702" => data <= "0001100111";
                when x"1703" => data <= "1111010110";
                when x"1704" => data <= "0001100111";
                when x"1705" => data <= "0101000100";
                when x"1706" => data <= "1100110111";
                when x"1707" => data <= "1111010110";
                when x"1708" => data <= "1111010110";
                when x"1709" => data <= "1111010110";
                when x"170A" => data <= "1011000000";
                when x"170B" => data <= "0101000100";
                when x"170C" => data <= "1011000000";
                when x"170D" => data <= "1000010100";
                when x"170E" => data <= "1010001000";
                when x"170F" => data <= "1010001000";
                when x"1710" => data <= "0001000101";
                when x"1711" => data <= "1010001000";
                when x"1712" => data <= "1010001000";
                when x"1713" => data <= "1101111111";
                when x"1714" => data <= "1101111111";
                when x"1715" => data <= "1101111111";
                when x"1716" => data <= "1101111111";
                when x"1717" => data <= "1101111111";
                when x"1718" => data <= "1110011110";
                when x"1719" => data <= "1011010111";
                when x"171A" => data <= "1010111101";
                when x"171B" => data <= "0011111011";
                when x"171C" => data <= "1101111111";
                when x"171D" => data <= "1101111111";
                when x"171E" => data <= "1101111111";
                when x"171F" => data <= "1010111101";
                when x"1720" => data <= "1101111111";
                when x"1721" => data <= "0100001100";
                when x"1722" => data <= "1101111111";
                when x"1723" => data <= "1101111111";
                when x"1724" => data <= "1000110110";
                when x"1725" => data <= "1101111111";
                when x"1726" => data <= "1011010111";
                when x"1727" => data <= "0001000101";
                when x"1728" => data <= "1101111111";
                when x"1729" => data <= "0001000101";
                when x"172A" => data <= "1101111111";
                when x"172B" => data <= "1010001000";
                when x"172C" => data <= "0110000111";
                when x"172D" => data <= "1011100010";
                when x"172E" => data <= "1100010101";
                when x"172F" => data <= "1101111111";
                when x"1730" => data <= "1101111111";
                when x"1731" => data <= "1101111111";
                when x"1732" => data <= "1101111111";
                when x"1733" => data <= "0000101111";
                when x"1734" => data <= "1101111111";
                when x"1735" => data <= "0100001100";
                when x"1736" => data <= "0011111011";
                when x"1737" => data <= "1010001000";
                when x"1738" => data <= "1101111111";
                when x"1739" => data <= "1010001000";
                when x"173A" => data <= "1101111111";
                when x"173B" => data <= "1101111111";
                when x"173C" => data <= "1101111111";
                when x"173D" => data <= "0110000111";
                when x"173E" => data <= "1101111111";
                when x"173F" => data <= "0100001100";
                when x"1740" => data <= "0001000101";
                when x"1741" => data <= "0011111011";
                when x"1742" => data <= "1101111111";
                when x"1743" => data <= "1101111111";
                when x"1744" => data <= "1101111111";
                when x"1745" => data <= "1101111111";
                when x"1746" => data <= "0111101101";
                when x"1747" => data <= "1101111111";
                when x"1748" => data <= "0111011000";
                when x"1749" => data <= "1010001000";
                when x"174A" => data <= "1011010111";
                when x"174B" => data <= "0111101101";
                when x"174C" => data <= "1010001000";
                when x"174D" => data <= "1010001000";
                when x"174E" => data <= "1100010101";
                when x"174F" => data <= "1101111111";
                when x"1750" => data <= "1010001000";
                when x"1751" => data <= "1101111111";
                when x"1752" => data <= "1010001000";
                when x"1753" => data <= "0000101111";
                when x"1754" => data <= "1101111111";
                when x"1755" => data <= "1101111111";
                when x"1756" => data <= "1101111111";
                when x"1757" => data <= "1010001000";
                when x"1758" => data <= "0011111011";
                when x"1759" => data <= "1101111111";
                when x"175A" => data <= "1010001000";
                when x"175B" => data <= "1010111101";
                when x"175C" => data <= "0000000000";
                when x"175D" => data <= "0000000000";
                when x"175E" => data <= "0000000000";
                when x"175F" => data <= "0000000000";
                when x"1760" => data <= "0000000000";
                when x"1761" => data <= "0000000000";
                when x"1762" => data <= "0000000000";
                when x"1763" => data <= "0000000000";
                when x"1764" => data <= "0000000000";
                when x"1765" => data <= "0000000000";
                when x"1766" => data <= "0000000000";
                when x"1767" => data <= "0000000000";
                when x"1768" => data <= "0000000000";
                when x"1769" => data <= "0000000000";
                when x"176A" => data <= "0000000000";
                when x"176B" => data <= "0000000000";
                when x"176C" => data <= "0000000000";
                when x"176D" => data <= "0000000000";
                when x"176E" => data <= "0000000000";
                when x"176F" => data <= "0000000000";
                when x"1770" => data <= "0000000000";
                when x"1771" => data <= "0000000000";
                when x"1772" => data <= "0000000000";
                when x"1773" => data <= "0000000000";
                when x"1774" => data <= "0000000000";
                when x"1775" => data <= "0000000000";
                when x"1776" => data <= "0000000000";
                when x"1777" => data <= "0000000000";
                when x"1778" => data <= "0000000000";
                when x"1779" => data <= "0000000000";
                when x"177A" => data <= "0000000000";
                when x"177B" => data <= "0000000000";
                when x"177C" => data <= "0000000000";
                when x"177D" => data <= "0000000000";
                when x"177E" => data <= "0000000000";
                when x"177F" => data <= "0000000000";
                when x"1780" => data <= "0000000000";
                when x"1781" => data <= "0000000000";
                when x"1782" => data <= "0000000000";
                when x"1783" => data <= "0000000000";
                when x"1784" => data <= "0000000000";
                when x"1785" => data <= "0000000000";
                when x"1786" => data <= "0000000000";
                when x"1787" => data <= "1111011011";
                when x"1788" => data <= "0000000000";
                when x"1789" => data <= "0000000000";
                when x"178A" => data <= "0000000000";
                when x"178B" => data <= "0000000000";
                when x"178C" => data <= "0000000000";
                when x"178D" => data <= "0000000000";
                when x"178E" => data <= "0000000000";
                when x"178F" => data <= "0000000000";
                when x"1790" => data <= "0000000000";
                when x"1791" => data <= "0000000000";
                when x"1792" => data <= "0000000000";
                when x"1793" => data <= "0000000000";
                when x"1794" => data <= "0000000000";
                when x"1795" => data <= "0000000000";
                when x"1796" => data <= "0000000000";
                when x"1797" => data <= "0000000000";
                when x"1798" => data <= "0000000000";
                when x"1799" => data <= "0000000000";
                when x"179A" => data <= "0000000000";
                when x"179B" => data <= "0000000000";
                when x"179C" => data <= "0000000000";
                when x"179D" => data <= "0111110111";
                when x"179E" => data <= "0000000000";
                when x"179F" => data <= "0000000000";
                when x"17A0" => data <= "0000000000";
                when x"17A1" => data <= "0000000000";
                when x"17A2" => data <= "0000000000";
                when x"17A3" => data <= "0000000000";
                when x"17A4" => data <= "0000000000";
                when x"17A5" => data <= "0000000000";
                when x"17A6" => data <= "0000000000";
                when x"17A7" => data <= "0000000000";
                when x"17A8" => data <= "0000000000";
                when x"17A9" => data <= "0000000000";
                when x"17AA" => data <= "0000000000";
                when x"17AB" => data <= "0000000000";
                when x"17AC" => data <= "0000000000";
                when x"17AD" => data <= "0000000000";
                when x"17AE" => data <= "0000000000";
                when x"17AF" => data <= "0000000000";
                when x"17B0" => data <= "0000000000";
                when x"17B1" => data <= "0000000000";
                when x"17B2" => data <= "0000000000";
                when x"17B3" => data <= "0000000000";
                when x"17B4" => data <= "0000000000";
                when x"17B5" => data <= "0000000000";
                when x"17B6" => data <= "0000000000";
                when x"17B7" => data <= "0000000000";
                when x"17B8" => data <= "0000000000";
                when x"17B9" => data <= "0000000000";
                when x"17BA" => data <= "0000000000";
                when x"17BB" => data <= "0000000000";
                when x"17BC" => data <= "0000000000";
                when x"17BD" => data <= "0000000000";
                when x"17BE" => data <= "0000000000";
                when x"17BF" => data <= "0000000000";
                when x"17C0" => data <= "0000000000";
                when x"17C1" => data <= "0000000000";
                when x"17C2" => data <= "0000000000";
                when x"17C3" => data <= "0000000000";
                when x"17C4" => data <= "0000000000";
                when x"17C5" => data <= "0000000000";
                when x"17C6" => data <= "0000000000";
                when x"17C7" => data <= "0000000000";
                when x"17C8" => data <= "0000000000";
                when x"17C9" => data <= "0000000000";
                when x"17CA" => data <= "0000000000";
                when x"17CB" => data <= "0000000000";
                when x"17CC" => data <= "0000000000";
                when x"17CD" => data <= "0000000000";
                when x"17CE" => data <= "0000000000";
                when x"17CF" => data <= "0000000000";
                when x"17D0" => data <= "0000000000";
                when x"17D1" => data <= "0000000000";
                when x"17D2" => data <= "0000000000";
                when x"17D3" => data <= "0000000000";
                when x"17D4" => data <= "0000000000";
                when x"17D5" => data <= "0000000000";
                when x"17D6" => data <= "0000000000";
                when x"17D7" => data <= "0000000000";
                when x"17D8" => data <= "0000000000";
                when x"17D9" => data <= "0000000000";
                when x"17DA" => data <= "0000000000";
                when x"17DB" => data <= "0000000000";
                when x"17DC" => data <= "0000000000";
                when x"17DD" => data <= "0000000000";
                when x"17DE" => data <= "0000000000";
                when x"17DF" => data <= "0000000000";
                when x"17E0" => data <= "1011001101";
                when x"17E1" => data <= "0000000000";
                when x"17E2" => data <= "0000000000";
                when x"17E3" => data <= "0000000000";
                when x"17E4" => data <= "0000000000";
                when x"17E5" => data <= "0000000000";
                when x"17E6" => data <= "0000000000";
                when x"17E7" => data <= "0000000000";
                when x"17E8" => data <= "0000000000";
                when x"17E9" => data <= "0000000000";
                when x"17EA" => data <= "0000000000";
                when x"17EB" => data <= "0000000000";
                when x"17EC" => data <= "0000000000";
                when x"17ED" => data <= "0000000000";
                when x"17EE" => data <= "0000000000";
                when x"17EF" => data <= "0000000000";
                when x"17F0" => data <= "0000000000";
                when x"17F1" => data <= "0000000000";
                when x"17F2" => data <= "0000000000";
                when x"17F3" => data <= "0000000000";
                when x"17F4" => data <= "0000000000";
                when x"17F5" => data <= "0000000000";
                when x"17F6" => data <= "0000000000";
                when x"17F7" => data <= "0000000000";
                when x"17F8" => data <= "0000000000";
                when x"17F9" => data <= "0000000000";
                when x"17FA" => data <= "0000000000";
                when x"17FB" => data <= "0000000000";
                when x"17FC" => data <= "0000000000";
                when x"17FD" => data <= "0000000000";
                when x"17FE" => data <= "0000000000";
                when x"17FF" => data <= "0000000000";
                when x"1800" => data <= "0000000000";
                when x"1801" => data <= "0000000000";
                when x"1802" => data <= "0000000000";
                when x"1803" => data <= "0000000000";
                when x"1804" => data <= "0000000000";
                when x"1805" => data <= "0000000000";
                when x"1806" => data <= "0000000000";
                when x"1807" => data <= "0000000000";
                when x"1808" => data <= "0000000000";
                when x"1809" => data <= "0000000000";
                when x"180A" => data <= "0000000000";
                when x"180B" => data <= "0000000000";
                when x"180C" => data <= "0000000000";
                when x"180D" => data <= "0000000000";
                when x"180E" => data <= "0000000000";
                when x"180F" => data <= "0000000000";
                when x"1810" => data <= "0000000000";
                when x"1811" => data <= "0000000000";
                when x"1812" => data <= "0000000000";
                when x"1813" => data <= "0000000000";
                when x"1814" => data <= "0000000000";
                when x"1815" => data <= "0000000000";
                when x"1816" => data <= "0000000000";
                when x"1817" => data <= "0000000000";
                when x"1818" => data <= "0000000000";
                when x"1819" => data <= "0000000000";
                when x"181A" => data <= "0000000000";
                when x"181B" => data <= "0000000000";
                when x"181C" => data <= "0000000000";
                when x"181D" => data <= "0000000000";
                when x"181E" => data <= "0000000000";
                when x"181F" => data <= "0000000000";
                when x"1820" => data <= "0000000000";
                when x"1821" => data <= "0000000000";
                when x"1822" => data <= "0000000000";
                when x"1823" => data <= "0000000000";
                when x"1824" => data <= "0000000000";
                when x"1825" => data <= "0000000000";
                when x"1826" => data <= "0000000000";
                when x"1827" => data <= "0000000000";
                when x"1828" => data <= "0000000000";
                when x"1829" => data <= "0000000000";
                when x"182A" => data <= "0000000000";
                when x"182B" => data <= "0000000000";
                when x"182C" => data <= "0000000000";
                when x"182D" => data <= "0000000000";
                when x"182E" => data <= "0000000000";
                when x"182F" => data <= "0000000000";
                when x"1830" => data <= "0000000000";
                when x"1831" => data <= "0000000000";
                when x"1832" => data <= "0000000000";
                when x"1833" => data <= "0000000000";
                when x"1834" => data <= "0000000000";
                when x"1835" => data <= "0000000000";
                when x"1836" => data <= "0000000000";
                when x"1837" => data <= "0000000000";
                when x"1838" => data <= "0100010110";
                when x"1839" => data <= "0000000000";
                when x"183A" => data <= "0000000000";
                when x"183B" => data <= "0000000000";
                when x"183C" => data <= "0000000000";
                when x"183D" => data <= "0000000000";
                when x"183E" => data <= "0000000000";
                when x"183F" => data <= "0000000000";
                when x"1840" => data <= "0000000000";
                when x"1841" => data <= "0000000000";
                when x"1842" => data <= "0000000000";
                when x"1843" => data <= "0000000000";
                when x"1844" => data <= "0000000000";
                when x"1845" => data <= "0000000000";
                when x"1846" => data <= "0000000000";
                when x"1847" => data <= "0000000000";
                when x"1848" => data <= "0000000000";
                when x"1849" => data <= "0000000000";
                when x"184A" => data <= "0000000000";
                when x"184B" => data <= "0000000000";
                when x"184C" => data <= "0000000000";
                when x"184D" => data <= "0000000000";
                when x"184E" => data <= "0000000000";
                when x"184F" => data <= "0000000000";
                when x"1850" => data <= "0000000000";
                when x"1851" => data <= "0000000000";
                when x"1852" => data <= "0000000000";
                when x"1853" => data <= "0000000000";
                when x"1854" => data <= "0000000000";
                when x"1855" => data <= "0000000000";
                when x"1856" => data <= "0000000000";
                when x"1857" => data <= "0000000000";
                when x"1858" => data <= "0000000000";
                when x"1859" => data <= "0000000000";
                when x"185A" => data <= "0000000000";
                when x"185B" => data <= "0000000000";
                when x"185C" => data <= "0000000000";
                when x"185D" => data <= "0000000000";
                when x"185E" => data <= "0000000000";
                when x"185F" => data <= "0000000000";
                when x"1860" => data <= "0000000000";
                when x"1861" => data <= "0000000000";
                when x"1862" => data <= "0000000000";
                when x"1863" => data <= "0000000000";
                when x"1864" => data <= "0000000000";
                when x"1865" => data <= "0000000000";
                when x"1866" => data <= "0000000000";
                when x"1867" => data <= "0000000000";
                when x"1868" => data <= "0000000000";
                when x"1869" => data <= "0000000000";
                when x"186A" => data <= "0000000000";
                when x"186B" => data <= "0000000000";
                when x"186C" => data <= "0000000000";
                when x"186D" => data <= "0000000000";
                when x"186E" => data <= "0000000000";
                when x"186F" => data <= "0000000000";
                when x"1870" => data <= "0000000000";
                when x"1871" => data <= "0000000000";
                when x"1872" => data <= "0000000000";
                when x"1873" => data <= "0000000000";
                when x"1874" => data <= "0000000000";
                when x"1875" => data <= "0000000000";
                when x"1876" => data <= "0000000000";
                when x"1877" => data <= "0000000000";
                when x"1878" => data <= "0000000000";
                when x"1879" => data <= "0000000000";
                when x"187A" => data <= "0000000000";
                when x"187B" => data <= "0000000000";
                when x"187C" => data <= "0000000000";
                when x"187D" => data <= "0000000000";
                when x"187E" => data <= "0000000000";
                when x"187F" => data <= "0000000000";
                when x"1880" => data <= "0000000000";
                when x"1881" => data <= "0000000000";
                when x"1882" => data <= "0000000000";
                when x"1883" => data <= "0000000000";
                when x"1884" => data <= "0000000000";
                when x"1885" => data <= "0000000000";
                when x"1886" => data <= "0000000000";
                when x"1887" => data <= "0000000000";
                when x"1888" => data <= "0000000000";
                when x"1889" => data <= "0000000000";
                when x"188A" => data <= "0000000000";
                when x"188B" => data <= "0000000000";
                when x"188C" => data <= "0000000000";
                when x"188D" => data <= "0000000000";
                when x"188E" => data <= "0000000000";
                when x"188F" => data <= "0000000000";
                when x"1890" => data <= "0000000000";
                when x"1891" => data <= "0000000000";
                when x"1892" => data <= "0000000000";
                when x"1893" => data <= "0000000000";
                when x"1894" => data <= "0000000000";
                when x"1895" => data <= "0000000000";
                when x"1896" => data <= "0000000000";
                when x"1897" => data <= "0000000000";
                when x"1898" => data <= "0000000000";
                when x"1899" => data <= "0000000000";
                when x"189A" => data <= "0000000000";
                when x"189B" => data <= "0000000000";
                when x"189C" => data <= "0000000000";
                when x"189D" => data <= "0000000000";
                when x"189E" => data <= "0000000000";
                when x"189F" => data <= "0000000000";
                when x"18A0" => data <= "0000000000";
                when x"18A1" => data <= "0000000000";
                when x"18A2" => data <= "0000000000";
                when x"18A3" => data <= "0000000000";
                when x"18A4" => data <= "0000000000";
                when x"18A5" => data <= "0000000000";
                when x"18A6" => data <= "0000000000";
                when x"18A7" => data <= "0000000000";
                when x"18A8" => data <= "0000000000";
                when x"18A9" => data <= "0000000000";
                when x"18AA" => data <= "0000000000";
                when x"18AB" => data <= "0000000000";
                when x"18AC" => data <= "0000000000";
                when x"18AD" => data <= "0000000000";
                when x"18AE" => data <= "0000000000";
                when x"18AF" => data <= "0000000000";
                when x"18B0" => data <= "0000000000";
                when x"18B1" => data <= "0000000000";
                when x"18B2" => data <= "0000000000";
                when x"18B3" => data <= "0000000000";
                when x"18B4" => data <= "0000000000";
                when x"18B5" => data <= "0000000000";
                when x"18B6" => data <= "0000000000";
                when x"18B7" => data <= "0000000000";
                when x"18B8" => data <= "0000000000";
                when x"18B9" => data <= "0000000000";
                when x"18BA" => data <= "0000000000";
                when x"18BB" => data <= "0000000000";
                when x"18BC" => data <= "0000000000";
                when x"18BD" => data <= "0000000000";
                when x"18BE" => data <= "0000000000";
                when x"18BF" => data <= "0000000000";
                when x"18C0" => data <= "0000000000";
                when x"18C1" => data <= "0000000000";
                when x"18C2" => data <= "0000000000";
                when x"18C3" => data <= "0000000000";
                when x"18C4" => data <= "0000000000";
                when x"18C5" => data <= "0000000000";
                when x"18C6" => data <= "0000000000";
                when x"18C7" => data <= "0000000000";
                when x"18C8" => data <= "0000000000";
                when x"18C9" => data <= "0000000000";
                when x"18CA" => data <= "0000000000";
                when x"18CB" => data <= "0000000000";
                when x"18CC" => data <= "0000000000";
                when x"18CD" => data <= "0000000000";
                when x"18CE" => data <= "0000000000";
                when x"18CF" => data <= "0000000000";
                when x"18D0" => data <= "0000000000";
                when x"18D1" => data <= "0000000000";
                when x"18D2" => data <= "0000000000";
                when x"18D3" => data <= "0000000000";
                when x"18D4" => data <= "0000000000";
                when x"18D5" => data <= "0000000000";
                when x"18D6" => data <= "0000000000";
                when x"18D7" => data <= "0000000000";
                when x"18D8" => data <= "0000000000";
                when x"18D9" => data <= "0000000000";
                when x"18DA" => data <= "0000000000";
                when x"18DB" => data <= "0000000000";
                when x"18DC" => data <= "0000000000";
                when x"18DD" => data <= "0000000000";
                when x"18DE" => data <= "0000000000";
                when x"18DF" => data <= "0000000000";
                when x"18E0" => data <= "0000000000";
                when x"18E1" => data <= "0000000000";
                when x"18E2" => data <= "0000000000";
                when x"18E3" => data <= "0000000000";
                when x"18E4" => data <= "0000000000";
                when x"18E5" => data <= "0000000000";
                when x"18E6" => data <= "0000000000";
                when x"18E7" => data <= "0000000000";
                when x"18E8" => data <= "0000000000";
                when x"18E9" => data <= "0000000000";
                when x"18EA" => data <= "0000000000";
                when x"18EB" => data <= "0000000000";
                when x"18EC" => data <= "0000000000";
                when x"18ED" => data <= "0000000000";
                when x"18EE" => data <= "0000000000";
                when x"18EF" => data <= "0000000000";
                when x"18F0" => data <= "0000000000";
                when x"18F1" => data <= "0000000000";
                when x"18F2" => data <= "0000000000";
                when x"18F3" => data <= "0000000000";
                when x"18F4" => data <= "0000000000";
                when x"18F5" => data <= "0000000000";
                when x"18F6" => data <= "0000000000";
                when x"18F7" => data <= "0000000000";
                when x"18F8" => data <= "0000000000";
                when x"18F9" => data <= "0000000000";
                when x"18FA" => data <= "0000000000";
                when x"18FB" => data <= "0000000000";
                when x"18FC" => data <= "0000000000";
                when x"18FD" => data <= "0000000000";
                when x"18FE" => data <= "0000000000";
                when x"18FF" => data <= "0000000000";
                when x"1900" => data <= "0000000000";
                when x"1901" => data <= "0000000000";
                when x"1902" => data <= "0000000000";
                when x"1903" => data <= "0000000000";
                when x"1904" => data <= "0000000000";
                when x"1905" => data <= "0000000000";
                when x"1906" => data <= "0000000000";
                when x"1907" => data <= "0000000000";
                when x"1908" => data <= "0000000000";
                when x"1909" => data <= "0000000000";
                when x"190A" => data <= "0000000000";
                when x"190B" => data <= "0000000000";
                when x"190C" => data <= "0000000000";
                when x"190D" => data <= "0000000000";
                when x"190E" => data <= "0000000000";
                when x"190F" => data <= "0000000000";
                when x"1910" => data <= "0000000000";
                when x"1911" => data <= "0000000000";
                when x"1912" => data <= "0000000000";
                when x"1913" => data <= "0000000000";
                when x"1914" => data <= "0000000000";
                when x"1915" => data <= "0000000000";
                when x"1916" => data <= "0000000000";
                when x"1917" => data <= "0000000000";
                when x"1918" => data <= "0000000000";
                when x"1919" => data <= "0000000000";
                when x"191A" => data <= "0000000000";
                when x"191B" => data <= "0000000000";
                when x"191C" => data <= "0000000000";
                when x"191D" => data <= "0000000000";
                when x"191E" => data <= "0000000000";
                when x"191F" => data <= "0000000000";
                when x"1920" => data <= "0000000000";
                when x"1921" => data <= "0000000000";
                when x"1922" => data <= "0000000000";
                when x"1923" => data <= "0000000000";
                when x"1924" => data <= "0000000000";
                when x"1925" => data <= "0000000000";
                when x"1926" => data <= "0111110111";
                when x"1927" => data <= "0000000000";
                when x"1928" => data <= "0000000000";
                when x"1929" => data <= "0000000000";
                when x"192A" => data <= "0000000000";
                when x"192B" => data <= "0000000000";
                when x"192C" => data <= "0000000000";
                when x"192D" => data <= "0000000000";
                when x"192E" => data <= "0000000000";
                when x"192F" => data <= "0000000000";
                when x"1930" => data <= "0000000000";
                when x"1931" => data <= "0000000000";
                when x"1932" => data <= "0000000000";
                when x"1933" => data <= "0000000000";
                when x"1934" => data <= "0000000000";
                when x"1935" => data <= "0000000000";
                when x"1936" => data <= "0000000000";
                when x"1937" => data <= "0000000000";
                when x"1938" => data <= "0000000000";
                when x"1939" => data <= "0000000000";
                when x"193A" => data <= "0000000000";
                when x"193B" => data <= "0000000000";
                when x"193C" => data <= "0000000000";
                when x"193D" => data <= "0000000000";
                when x"193E" => data <= "0000000000";
                when x"193F" => data <= "0000000000";
                when x"1940" => data <= "0000000000";
                when x"1941" => data <= "0000000000";
                when x"1942" => data <= "0000000000";
                when x"1943" => data <= "0000000000";
                when x"1944" => data <= "0000000000";
                when x"1945" => data <= "0000000000";
                when x"1946" => data <= "0000000000";
                when x"1947" => data <= "0000000000";
                when x"1948" => data <= "0000000000";
                when x"1949" => data <= "0000000000";
                when x"194A" => data <= "0000000000";
                when x"194B" => data <= "0000000000";
                when x"194C" => data <= "0000000000";
                when x"194D" => data <= "0000000000";
                when x"194E" => data <= "0000000000";
                when x"194F" => data <= "0000000000";
                when x"1950" => data <= "0000000000";
                when x"1951" => data <= "0000000000";
                when x"1952" => data <= "0000000000";
                when x"1953" => data <= "0000000000";
                when x"1954" => data <= "0000000000";
                when x"1955" => data <= "0000000000";
                when x"1956" => data <= "0000000000";
                when x"1957" => data <= "0000000000";
                when x"1958" => data <= "0000000000";
                when x"1959" => data <= "0000000000";
                when x"195A" => data <= "0000000000";
                when x"195B" => data <= "0000000000";
                when x"195C" => data <= "0000000000";
                when x"195D" => data <= "0000000000";
                when x"195E" => data <= "0000000000";
                when x"195F" => data <= "0000000000";
                when x"1960" => data <= "0000000000";
                when x"1961" => data <= "0000000000";
                when x"1962" => data <= "0000000000";
                when x"1963" => data <= "0000000000";
                when x"1964" => data <= "0000000000";
                when x"1965" => data <= "0000000000";
                when x"1966" => data <= "0000000000";
                when x"1967" => data <= "0000000000";
                when x"1968" => data <= "0000000000";
                when x"1969" => data <= "0000000000";
                when x"196A" => data <= "0000000000";
                when x"196B" => data <= "0000000000";
                when x"196C" => data <= "0000000000";
                when x"196D" => data <= "0000000000";
                when x"196E" => data <= "0000000000";
                when x"196F" => data <= "0000000000";
                when x"1970" => data <= "0000000000";
                when x"1971" => data <= "0000000000";
                when x"1972" => data <= "0000000000";
                when x"1973" => data <= "0000000000";
                when x"1974" => data <= "0000000000";
                when x"1975" => data <= "0000000000";
                when x"1976" => data <= "0000000000";
                when x"1977" => data <= "0000000000";
                when x"1978" => data <= "0000000000";
                when x"1979" => data <= "0000000000";
                when x"197A" => data <= "0000000000";
                when x"197B" => data <= "0000000000";
                when x"197C" => data <= "0000000000";
                when x"197D" => data <= "0000000000";
                when x"197E" => data <= "0000000000";
                when x"197F" => data <= "0000000000";
                when x"1980" => data <= "0000000000";
                when x"1981" => data <= "0000000000";
                when x"1982" => data <= "0000000000";
                when x"1983" => data <= "0000000000";
                when x"1984" => data <= "0000000000";
                when x"1985" => data <= "0000000000";
                when x"1986" => data <= "0000000000";
                when x"1987" => data <= "0000000000";
                when x"1988" => data <= "0000000000";
                when x"1989" => data <= "0000000000";
                when x"198A" => data <= "0000000000";
                when x"198B" => data <= "0000000000";
                when x"198C" => data <= "0000000000";
                when x"198D" => data <= "0000000000";
                when x"198E" => data <= "0000000000";
                when x"198F" => data <= "0000000000";
                when x"1990" => data <= "0000000000";
                when x"1991" => data <= "0000000000";
                when x"1992" => data <= "0000000000";
                when x"1993" => data <= "0000000000";
                when x"1994" => data <= "0000000000";
                when x"1995" => data <= "0000000000";
                when x"1996" => data <= "0000000000";
                when x"1997" => data <= "0000000000";
                when x"1998" => data <= "0000000000";
                when x"1999" => data <= "0000000000";
                when x"199A" => data <= "0000000000";
                when x"199B" => data <= "0000000000";
                when x"199C" => data <= "0000000000";
                when x"199D" => data <= "0000000000";
                when x"199E" => data <= "0000000000";
                when x"199F" => data <= "0000000000";
                when x"19A0" => data <= "0000000000";
                when x"19A1" => data <= "0000000000";
                when x"19A2" => data <= "0000000000";
                when x"19A3" => data <= "0000000000";
                when x"19A4" => data <= "0000000000";
                when x"19A5" => data <= "0000000000";
                when x"19A6" => data <= "0000000000";
                when x"19A7" => data <= "0000000000";
                when x"19A8" => data <= "0000000000";
                when x"19A9" => data <= "0000000000";
                when x"19AA" => data <= "0000000000";
                when x"19AB" => data <= "0000000000";
                when x"19AC" => data <= "0000000000";
                when x"19AD" => data <= "0000000000";
                when x"19AE" => data <= "0000000000";
                when x"19AF" => data <= "0000000000";
                when x"19B0" => data <= "0000000000";
                when x"19B1" => data <= "0000000000";
                when x"19B2" => data <= "0000000000";
                when x"19B3" => data <= "0000000000";
                when x"19B4" => data <= "0000000000";
                when x"19B5" => data <= "0000000000";
                when x"19B6" => data <= "0000000000";
                when x"19B7" => data <= "0000000000";
                when x"19B8" => data <= "0000000000";
                when x"19B9" => data <= "0000000000";
                when x"19BA" => data <= "0000000000";
                when x"19BB" => data <= "0000000000";
                when x"19BC" => data <= "0000000000";
                when x"19BD" => data <= "0000000000";
                when x"19BE" => data <= "0000000000";
                when x"19BF" => data <= "0000000000";
                when x"19C0" => data <= "0000000000";
                when x"19C1" => data <= "0000000000";
                when x"19C2" => data <= "0000000000";
                when x"19C3" => data <= "0000000000";
                when x"19C4" => data <= "0000000000";
                when x"19C5" => data <= "0000000000";
                when x"19C6" => data <= "0000000000";
                when x"19C7" => data <= "0000000000";
                when x"19C8" => data <= "0000000000";
                when x"19C9" => data <= "0000000000";
                when x"19CA" => data <= "0000000000";
                when x"19CB" => data <= "0000000000";
                when x"19CC" => data <= "0000000000";
                when x"19CD" => data <= "0000000000";
                when x"19CE" => data <= "0000000000";
                when x"19CF" => data <= "0000000000";
                when x"19D0" => data <= "0000000000";
                when x"19D1" => data <= "0000000000";
                when x"19D2" => data <= "0000000000";
                when x"19D3" => data <= "0000000000";
                when x"19D4" => data <= "0000000000";
                when x"19D5" => data <= "0000000000";
                when x"19D6" => data <= "0000000000";
                when x"19D7" => data <= "0000000000";
                when x"19D8" => data <= "0000000000";
                when x"19D9" => data <= "0000000000";
                when x"19DA" => data <= "0000000000";
                when x"19DB" => data <= "0000000000";
                when x"19DC" => data <= "0000000000";
                when x"19DD" => data <= "0000000000";
                when x"19DE" => data <= "0000000000";
                when x"19DF" => data <= "0000000000";
                when x"19E0" => data <= "0000000000";
                when x"19E1" => data <= "0000000000";
                when x"19E2" => data <= "0000000000";
                when x"19E3" => data <= "0000000000";
                when x"19E4" => data <= "0000000000";
                when x"19E5" => data <= "0000000000";
                when x"19E6" => data <= "0000000000";
                when x"19E7" => data <= "0000000000";
                when x"19E8" => data <= "0000000000";
                when x"19E9" => data <= "0000000000";
                when x"19EA" => data <= "0000000000";
                when x"19EB" => data <= "0000000000";
                when x"19EC" => data <= "0000000000";
                when x"19ED" => data <= "0000000000";
                when x"19EE" => data <= "0000000000";
                when x"19EF" => data <= "0000000000";
                when x"19F0" => data <= "0000000000";
                when x"19F1" => data <= "0000000000";
                when x"19F2" => data <= "0000000000";
                when x"19F3" => data <= "0000000000";
                when x"19F4" => data <= "0000000000";
                when x"19F5" => data <= "0000000000";
                when x"19F6" => data <= "0000000000";
                when x"19F7" => data <= "0000000000";
                when x"19F8" => data <= "0000000000";
                when x"19F9" => data <= "0000000000";
                when x"19FA" => data <= "0000000000";
                when x"19FB" => data <= "0000000000";
                when x"19FC" => data <= "0000000000";
                when x"19FD" => data <= "0000000000";
                when x"19FE" => data <= "0000000000";
                when x"19FF" => data <= "0000000000";
                when x"1A00" => data <= "0000000000";
                when x"1A01" => data <= "0000000000";
                when x"1A02" => data <= "0000000000";
                when x"1A03" => data <= "0000000000";
                when x"1A04" => data <= "0000000000";
                when x"1A05" => data <= "0000000000";
                when x"1A06" => data <= "0000000000";
                when x"1A07" => data <= "0000000000";
                when x"1A08" => data <= "0000000000";
                when x"1A09" => data <= "0000000000";
                when x"1A0A" => data <= "0000000000";
                when x"1A0B" => data <= "0000000000";
                when x"1A0C" => data <= "0000000000";
                when x"1A0D" => data <= "0000000000";
                when x"1A0E" => data <= "0000000000";
                when x"1A0F" => data <= "0000000000";
                when x"1A10" => data <= "0000000000";
                when x"1A11" => data <= "0000000000";
                when x"1A12" => data <= "0000000000";
                when x"1A13" => data <= "0000000000";
                when x"1A14" => data <= "0000000000";
                when x"1A15" => data <= "0000000000";
                when x"1A16" => data <= "0000000000";
                when x"1A17" => data <= "0000000000";
                when x"1A18" => data <= "0000000000";
                when x"1A19" => data <= "0000000000";
                when x"1A1A" => data <= "0000000000";
                when x"1A1B" => data <= "0000000000";
                when x"1A1C" => data <= "0000000000";
                when x"1A1D" => data <= "0000000000";
                when x"1A1E" => data <= "0000000000";
                when x"1A1F" => data <= "0000000000";
                when x"1A20" => data <= "0000000000";
                when x"1A21" => data <= "0000000000";
                when x"1A22" => data <= "0000000000";
                when x"1A23" => data <= "0000000000";
                when x"1A24" => data <= "0000000000";
                when x"1A25" => data <= "0000000000";
                when x"1A26" => data <= "0000000000";
                when x"1A27" => data <= "0000000000";
                when x"1A28" => data <= "0000000000";
                when x"1A29" => data <= "0000000000";
                when x"1A2A" => data <= "0000000000";
                when x"1A2B" => data <= "0000000000";
                when x"1A2C" => data <= "0000000000";
                when x"1A2D" => data <= "0000000000";
                when x"1A2E" => data <= "0000000000";
                when x"1A2F" => data <= "0000000000";
                when x"1A30" => data <= "0000000000";
                when x"1A31" => data <= "0000000000";
                when x"1A32" => data <= "0000000000";
                when x"1A33" => data <= "0000000000";
                when x"1A34" => data <= "0000000000";
                when x"1A35" => data <= "0000000000";
                when x"1A36" => data <= "0000000000";
                when x"1A37" => data <= "0000000000";
                when x"1A38" => data <= "0000000000";
                when x"1A39" => data <= "0000000000";
                when x"1A3A" => data <= "0000000000";
                when x"1A3B" => data <= "0000000000";
                when x"1A3C" => data <= "0000000000";
                when x"1A3D" => data <= "0000000000";
                when x"1A3E" => data <= "0000000000";
                when x"1A3F" => data <= "0000000000";
                when x"1A40" => data <= "0000000000";
                when x"1A41" => data <= "0000000000";
                when x"1A42" => data <= "0000000000";
                when x"1A43" => data <= "0000000000";
                when x"1A44" => data <= "0000000000";
                when x"1A45" => data <= "0000000000";
                when x"1A46" => data <= "0000000000";
                when x"1A47" => data <= "0000000000";
                when x"1A48" => data <= "0000000000";
                when x"1A49" => data <= "0000000000";
                when x"1A4A" => data <= "0000000000";
                when x"1A4B" => data <= "0000000000";
                when x"1A4C" => data <= "0000000000";
                when x"1A4D" => data <= "0000000000";
                when x"1A4E" => data <= "0000000000";
                when x"1A4F" => data <= "0000000000";
                when x"1A50" => data <= "0000000000";
                when x"1A51" => data <= "0000000000";
                when x"1A52" => data <= "0000000000";
                when x"1A53" => data <= "0000000000";
                when x"1A54" => data <= "0000000000";
                when x"1A55" => data <= "0000000000";
                when x"1A56" => data <= "0000000000";
                when x"1A57" => data <= "0000000000";
                when x"1A58" => data <= "0000000000";
                when x"1A59" => data <= "0000000000";
                when x"1A5A" => data <= "0000000000";
                when x"1A5B" => data <= "0000000000";
                when x"1A5C" => data <= "0000000000";
                when x"1A5D" => data <= "0000000000";
                when x"1A5E" => data <= "0000000000";
                when x"1A5F" => data <= "0000000000";
                when x"1A60" => data <= "0000000000";
                when x"1A61" => data <= "0000000000";
                when x"1A62" => data <= "0000000000";
                when x"1A63" => data <= "0000000000";
                when x"1A64" => data <= "0000000000";
                when x"1A65" => data <= "0000000000";
                when x"1A66" => data <= "0000000000";
                when x"1A67" => data <= "0000000000";
                when x"1A68" => data <= "0000000000";
                when x"1A69" => data <= "0000000000";
                when x"1A6A" => data <= "0000000000";
                when x"1A6B" => data <= "0000000000";
                when x"1A6C" => data <= "0000000000";
                when x"1A6D" => data <= "0000000000";
                when x"1A6E" => data <= "0000000000";
                when x"1A6F" => data <= "0000000000";
                when x"1A70" => data <= "0000000000";
                when x"1A71" => data <= "0000000000";
                when x"1A72" => data <= "0000000000";
                when x"1A73" => data <= "0000000000";
                when x"1A74" => data <= "0000000000";
                when x"1A75" => data <= "0000000000";
                when x"1A76" => data <= "0000000000";
                when x"1A77" => data <= "0000000000";
                when x"1A78" => data <= "0000000000";
                when x"1A79" => data <= "0000000000";
                when x"1A7A" => data <= "0000000000";
                when x"1A7B" => data <= "0000000000";
                when x"1A7C" => data <= "0000000000";
                when x"1A7D" => data <= "0000000000";
                when x"1A7E" => data <= "0000000000";
                when x"1A7F" => data <= "0000000000";
                when x"1A80" => data <= "0000000000";
                when x"1A81" => data <= "0000000000";
                when x"1A82" => data <= "0000000000";
                when x"1A83" => data <= "0000000000";
                when x"1A84" => data <= "0000000000";
                when x"1A85" => data <= "0000000000";
                when x"1A86" => data <= "0000000000";
                when x"1A87" => data <= "0000000000";
                when x"1A88" => data <= "0000000000";
                when x"1A89" => data <= "0000000000";
                when x"1A8A" => data <= "0000000000";
                when x"1A8B" => data <= "0000000000";
                when x"1A8C" => data <= "0000000000";
                when x"1A8D" => data <= "0000000000";
                when x"1A8E" => data <= "0000000000";
                when x"1A8F" => data <= "0000000000";
                when x"1A90" => data <= "0000000000";
                when x"1A91" => data <= "0000000000";
                when x"1A92" => data <= "0000000000";
                when x"1A93" => data <= "0000000000";
                when x"1A94" => data <= "0000000000";
                when x"1A95" => data <= "0000000000";
                when x"1A96" => data <= "0000000000";
                when x"1A97" => data <= "0000000000";
                when x"1A98" => data <= "0000000000";
                when x"1A99" => data <= "0000000000";
                when x"1A9A" => data <= "0000000000";
                when x"1A9B" => data <= "0000000000";
                when x"1A9C" => data <= "0000000000";
                when x"1A9D" => data <= "0000000000";
                when x"1A9E" => data <= "0000000000";
                when x"1A9F" => data <= "0000000000";
                when x"1AA0" => data <= "0000000000";
                when x"1AA1" => data <= "0000000000";
                when x"1AA2" => data <= "0000000000";
                when x"1AA3" => data <= "0000000000";
                when x"1AA4" => data <= "0000000000";
                when x"1AA5" => data <= "0000000000";
                when x"1AA6" => data <= "0000000000";
                when x"1AA7" => data <= "0000000000";
                when x"1AA8" => data <= "0000000000";
                when x"1AA9" => data <= "0000000000";
                when x"1AAA" => data <= "0000000000";
                when x"1AAB" => data <= "0000000000";
                when x"1AAC" => data <= "0000000000";
                when x"1AAD" => data <= "0000000000";
                when x"1AAE" => data <= "0000000000";
                when x"1AAF" => data <= "0000000000";
                when x"1AB0" => data <= "0000000000";
                when x"1AB1" => data <= "0000000000";
                when x"1AB2" => data <= "0000000000";
                when x"1AB3" => data <= "0000000000";
                when x"1AB4" => data <= "0000000000";
                when x"1AB5" => data <= "0000000000";
                when x"1AB6" => data <= "0000000000";
                when x"1AB7" => data <= "0000000000";
                when x"1AB8" => data <= "0000000000";
                when x"1AB9" => data <= "0000000000";
                when x"1ABA" => data <= "0000000000";
                when x"1ABB" => data <= "0000000000";
                when x"1ABC" => data <= "0000000000";
                when x"1ABD" => data <= "0000000000";
                when x"1ABE" => data <= "0000000000";
                when x"1ABF" => data <= "0000000000";
                when x"1AC0" => data <= "0000000000";
                when x"1AC1" => data <= "0000000000";
                when x"1AC2" => data <= "0000000000";
                when x"1AC3" => data <= "0000000000";
                when x"1AC4" => data <= "0000000000";
                when x"1AC5" => data <= "0000000000";
                when x"1AC6" => data <= "0000000000";
                when x"1AC7" => data <= "0000000000";
                when x"1AC8" => data <= "0000000000";
                when x"1AC9" => data <= "0000000000";
                when x"1ACA" => data <= "0000000000";
                when x"1ACB" => data <= "0000000000";
                when x"1ACC" => data <= "0000000000";
                when x"1ACD" => data <= "0000000000";
                when x"1ACE" => data <= "0000000000";
                when x"1ACF" => data <= "0000000000";
                when x"1AD0" => data <= "0000000000";
                when x"1AD1" => data <= "0000000000";
                when x"1AD2" => data <= "0000000000";
                when x"1AD3" => data <= "0000000000";
                when x"1AD4" => data <= "0000000000";
                when x"1AD5" => data <= "0000000000";
                when x"1AD6" => data <= "0000000000";
                when x"1AD7" => data <= "0000000000";
                when x"1AD8" => data <= "0000000000";
                when x"1AD9" => data <= "0000000000";
                when x"1ADA" => data <= "0000000000";
                when x"1ADB" => data <= "0000000000";
                when x"1ADC" => data <= "0000000000";
                when x"1ADD" => data <= "0000000000";
                when x"1ADE" => data <= "0000000000";
                when x"1ADF" => data <= "0000000000";
                when x"1AE0" => data <= "0000000000";
                when x"1AE1" => data <= "0000000000";
                when x"1AE2" => data <= "0000000000";
                when x"1AE3" => data <= "0000000000";
                when x"1AE4" => data <= "0000000000";
                when x"1AE5" => data <= "0000000000";
                when x"1AE6" => data <= "0000000000";
                when x"1AE7" => data <= "0000000000";
                when x"1AE8" => data <= "0000000000";
                when x"1AE9" => data <= "0000000000";
                when x"1AEA" => data <= "0000000000";
                when x"1AEB" => data <= "0000000000";
                when x"1AEC" => data <= "0000000000";
                when x"1AED" => data <= "0000000000";
                when x"1AEE" => data <= "0111110111";
                when x"1AEF" => data <= "0000000000";
                when x"1AF0" => data <= "0000000000";
                when x"1AF1" => data <= "0000000000";
                when x"1AF2" => data <= "0000000000";
                when x"1AF3" => data <= "0000000000";
                when x"1AF4" => data <= "0000000000";
                when x"1AF5" => data <= "0000000000";
                when x"1AF6" => data <= "0000000000";
                when x"1AF7" => data <= "0000000000";
                when x"1AF8" => data <= "0000000000";
                when x"1AF9" => data <= "0000000000";
                when x"1AFA" => data <= "0000000000";
                when x"1AFB" => data <= "0000000000";
                when x"1AFC" => data <= "0000000000";
                when x"1AFD" => data <= "0000000000";
                when x"1AFE" => data <= "0000000000";
                when x"1AFF" => data <= "0000000000";
                when x"1B00" => data <= "0000000000";
                when x"1B01" => data <= "0000000000";
                when x"1B02" => data <= "0000000000";
                when x"1B03" => data <= "0000000000";
                when x"1B04" => data <= "0000000000";
                when x"1B05" => data <= "0000000000";
                when x"1B06" => data <= "0000000000";
                when x"1B07" => data <= "0000000000";
                when x"1B08" => data <= "0000000000";
                when x"1B09" => data <= "0000000000";
                when x"1B0A" => data <= "0000000000";
                when x"1B0B" => data <= "0000000000";
                when x"1B0C" => data <= "0000000000";
                when x"1B0D" => data <= "0000000000";
                when x"1B0E" => data <= "0000000000";
                when x"1B0F" => data <= "0000000000";
                when x"1B10" => data <= "0000000000";
                when x"1B11" => data <= "0000000000";
                when x"1B12" => data <= "0000000000";
                when x"1B13" => data <= "0000000000";
                when x"1B14" => data <= "0000000000";
                when x"1B15" => data <= "0000000000";
                when x"1B16" => data <= "0000000000";
                when x"1B17" => data <= "0000000000";
                when x"1B18" => data <= "0000000000";
                when x"1B19" => data <= "0000000000";
                when x"1B1A" => data <= "0000000000";
                when x"1B1B" => data <= "0000000000";
                when x"1B1C" => data <= "0000000000";
                when x"1B1D" => data <= "0000000000";
                when x"1B1E" => data <= "0000000000";
                when x"1B1F" => data <= "0000000000";
                when x"1B20" => data <= "0000000000";
                when x"1B21" => data <= "0000000000";
                when x"1B22" => data <= "0000000000";
                when x"1B23" => data <= "0000000000";
                when x"1B24" => data <= "0000000000";
                when x"1B25" => data <= "0000000000";
                when x"1B26" => data <= "0000000000";
                when x"1B27" => data <= "0000000000";
                when x"1B28" => data <= "0000000000";
                when x"1B29" => data <= "0000000000";
                when x"1B2A" => data <= "0000000000";
                when x"1B2B" => data <= "0000000000";
                when x"1B2C" => data <= "0000000000";
                when x"1B2D" => data <= "0000000000";
                when x"1B2E" => data <= "0000000000";
                when x"1B2F" => data <= "0000000000";
                when x"1B30" => data <= "0000000000";
                when x"1B31" => data <= "0000000000";
                when x"1B32" => data <= "0000000000";
                when x"1B33" => data <= "0000000000";
                when x"1B34" => data <= "0000000000";
                when x"1B35" => data <= "0000000000";
                when x"1B36" => data <= "0000000000";
                when x"1B37" => data <= "0000000000";
                when x"1B38" => data <= "0000000000";
                when x"1B39" => data <= "0000000000";
                when x"1B3A" => data <= "0000000000";
                when x"1B3B" => data <= "0000000000";
                when x"1B3C" => data <= "0000000000";
                when x"1B3D" => data <= "0000000000";
                when x"1B3E" => data <= "0000000000";
                when x"1B3F" => data <= "0000000000";
                when x"1B40" => data <= "0000000000";
                when x"1B41" => data <= "0000000000";
                when x"1B42" => data <= "0000000000";
                when x"1B43" => data <= "0000000000";
                when x"1B44" => data <= "0000000000";
                when x"1B45" => data <= "0000000000";
                when x"1B46" => data <= "0000000000";
                when x"1B47" => data <= "0000000000";
                when x"1B48" => data <= "0000000000";
                when x"1B49" => data <= "0000000000";
                when x"1B4A" => data <= "0000000000";
                when x"1B4B" => data <= "0000000000";
                when x"1B4C" => data <= "0000000000";
                when x"1B4D" => data <= "0000000000";
                when x"1B4E" => data <= "0000000000";
                when x"1B4F" => data <= "0000000000";
                when x"1B50" => data <= "0000000000";
                when x"1B51" => data <= "0000000000";
                when x"1B52" => data <= "0000000000";
                when x"1B53" => data <= "0000000000";
                when x"1B54" => data <= "0000000000";
                when x"1B55" => data <= "0000000000";
                when x"1B56" => data <= "0000000000";
                when x"1B57" => data <= "0000000000";
                when x"1B58" => data <= "0000000000";
                when x"1B59" => data <= "0000000000";
                when x"1B5A" => data <= "0000000000";
                when x"1B5B" => data <= "0000000000";
                when x"1B5C" => data <= "0000000000";
                when x"1B5D" => data <= "0000000000";
                when x"1B5E" => data <= "0000000000";
                when x"1B5F" => data <= "0000000000";
                when x"1B60" => data <= "0000000000";
                when x"1B61" => data <= "0000000000";
                when x"1B62" => data <= "0000000000";
                when x"1B63" => data <= "0000000000";
                when x"1B64" => data <= "0000000000";
                when x"1B65" => data <= "0000000000";
                when x"1B66" => data <= "0000000000";
                when x"1B67" => data <= "0000000000";
                when x"1B68" => data <= "0000000000";
                when x"1B69" => data <= "0000000000";
                when x"1B6A" => data <= "0000000000";
                when x"1B6B" => data <= "0000000000";
                when x"1B6C" => data <= "0000000000";
                when x"1B6D" => data <= "0000000000";
                when x"1B6E" => data <= "0000000000";
                when x"1B6F" => data <= "0000000000";
                when x"1B70" => data <= "0000000000";
                when x"1B71" => data <= "0000000000";
                when x"1B72" => data <= "0000000000";
                when x"1B73" => data <= "0000000000";
                when x"1B74" => data <= "0000000000";
                when x"1B75" => data <= "0000000000";
                when x"1B76" => data <= "0000000000";
                when x"1B77" => data <= "0000000000";
                when x"1B78" => data <= "0000000000";
                when x"1B79" => data <= "0000000000";
                when x"1B7A" => data <= "0000000000";
                when x"1B7B" => data <= "0000000000";
                when x"1B7C" => data <= "0000000000";
                when x"1B7D" => data <= "0000000000";
                when x"1B7E" => data <= "0000000000";
                when x"1B7F" => data <= "0000000000";
                when x"1B80" => data <= "0000000000";
                when x"1B81" => data <= "1010100111";
                when x"1B82" => data <= "0000000000";
                when x"1B83" => data <= "0000000000";
                when x"1B84" => data <= "0000000000";
                when x"1B85" => data <= "0000000000";
                when x"1B86" => data <= "0000000000";
                when x"1B87" => data <= "0000000000";
                when x"1B88" => data <= "0000000000";
                when x"1B89" => data <= "0000000000";
                when x"1B8A" => data <= "0000000000";
                when x"1B8B" => data <= "0000000000";
                when x"1B8C" => data <= "0000000000";
                when x"1B8D" => data <= "0000000000";
                when x"1B8E" => data <= "0000000000";
                when x"1B8F" => data <= "0000000000";
                when x"1B90" => data <= "0000000000";
                when x"1B91" => data <= "0000000000";
                when x"1B92" => data <= "0000000000";
                when x"1B93" => data <= "0000000000";
                when x"1B94" => data <= "0000000000";
                when x"1B95" => data <= "0000000000";
                when x"1B96" => data <= "0000000000";
                when x"1B97" => data <= "0000000000";
                when x"1B98" => data <= "0000000000";
                when x"1B99" => data <= "0000000000";
                when x"1B9A" => data <= "0000000000";
                when x"1B9B" => data <= "0000000000";
                when x"1B9C" => data <= "0000000000";
                when x"1B9D" => data <= "0000000000";
                when x"1B9E" => data <= "0000000000";
                when x"1B9F" => data <= "0000000000";
                when x"1BA0" => data <= "0000000000";
                when x"1BA1" => data <= "0000000000";
                when x"1BA2" => data <= "0000000000";
                when x"1BA3" => data <= "0000000000";
                when x"1BA4" => data <= "0000000000";
                when x"1BA5" => data <= "0000000000";
                when x"1BA6" => data <= "0000000000";
                when x"1BA7" => data <= "0000000000";
                when x"1BA8" => data <= "0000000000";
                when x"1BA9" => data <= "0000000000";
                when x"1BAA" => data <= "0000000000";
                when x"1BAB" => data <= "0000000000";
                when x"1BAC" => data <= "0000000000";
                when x"1BAD" => data <= "0000000000";
                when x"1BAE" => data <= "0000000000";
                when x"1BAF" => data <= "0000000000";
                when x"1BB0" => data <= "0000000000";
                when x"1BB1" => data <= "0000000000";
                when x"1BB2" => data <= "0000000000";
                when x"1BB3" => data <= "0000000000";
                when x"1BB4" => data <= "0000000000";
                when x"1BB5" => data <= "0000000000";
                when x"1BB6" => data <= "0000000000";
                when x"1BB7" => data <= "0000000000";
                when x"1BB8" => data <= "0000000000";
                when x"1BB9" => data <= "0000000000";
                when x"1BBA" => data <= "0000000000";
                when x"1BBB" => data <= "0000000000";
                when x"1BBC" => data <= "0000000000";
                when x"1BBD" => data <= "0000000000";
                when x"1BBE" => data <= "0000000000";
                when x"1BBF" => data <= "0000000000";
                when x"1BC0" => data <= "0000000000";
                when x"1BC1" => data <= "0000000000";
                when x"1BC2" => data <= "0000000000";
                when x"1BC3" => data <= "0000000000";
                when x"1BC4" => data <= "0000000000";
                when x"1BC5" => data <= "0000000000";
                when x"1BC6" => data <= "0000000000";
                when x"1BC7" => data <= "0000000000";
                when x"1BC8" => data <= "0000000000";
                when x"1BC9" => data <= "0000000000";
                when x"1BCA" => data <= "0000000000";
                when x"1BCB" => data <= "0000000000";
                when x"1BCC" => data <= "0000000000";
                when x"1BCD" => data <= "0000000000";
                when x"1BCE" => data <= "0000000000";
                when x"1BCF" => data <= "0000000000";
                when x"1BD0" => data <= "0000000000";
                when x"1BD1" => data <= "0000000000";
                when x"1BD2" => data <= "0000000000";
                when x"1BD3" => data <= "0000000000";
                when x"1BD4" => data <= "0000000000";
                when x"1BD5" => data <= "0000000000";
                when x"1BD6" => data <= "0000000000";
                when x"1BD7" => data <= "0000000000";
                when x"1BD8" => data <= "0000000000";
                when x"1BD9" => data <= "0000000000";
                when x"1BDA" => data <= "0000000000";
                when x"1BDB" => data <= "1011001101";
                when x"1BDC" => data <= "0000000000";
                when x"1BDD" => data <= "0000000000";
                when x"1BDE" => data <= "0000000000";
                when x"1BDF" => data <= "0000000000";
                when x"1BE0" => data <= "0000000000";
                when x"1BE1" => data <= "0000000000";
                when x"1BE2" => data <= "0000000000";
                when x"1BE3" => data <= "0000000000";
                when x"1BE4" => data <= "0000000000";
                when x"1BE5" => data <= "0000000000";
                when x"1BE6" => data <= "0000000000";
                when x"1BE7" => data <= "0000000000";
                when x"1BE8" => data <= "0000000000";
                when x"1BE9" => data <= "0000000000";
                when x"1BEA" => data <= "0000000000";
                when x"1BEB" => data <= "0000000000";
                when x"1BEC" => data <= "0000000000";
                when x"1BED" => data <= "0000000000";
                when x"1BEE" => data <= "0000000000";
                when x"1BEF" => data <= "0000000000";
                when x"1BF0" => data <= "0000000000";
                when x"1BF1" => data <= "0000000000";
                when x"1BF2" => data <= "0000000000";
                when x"1BF3" => data <= "0000000000";
                when x"1BF4" => data <= "0000000000";
                when x"1BF5" => data <= "0000000000";
                when x"1BF6" => data <= "0000000000";
                when x"1BF7" => data <= "0000000000";
                when x"1BF8" => data <= "0000000000";
                when x"1BF9" => data <= "0000000000";
                when x"1BFA" => data <= "0000000000";
                when x"1BFB" => data <= "0000000000";
                when x"1BFC" => data <= "0000000000";
                when x"1BFD" => data <= "0000000000";
                when x"1BFE" => data <= "0000000000";
                when x"1BFF" => data <= "0000000000";
                when x"1C00" => data <= "0000000000";
                when x"1C01" => data <= "0000000000";
                when x"1C02" => data <= "0000000000";
                when x"1C03" => data <= "0000000000";
                when x"1C04" => data <= "0000000000";
                when x"1C05" => data <= "0000000000";
                when x"1C06" => data <= "0000000000";
                when x"1C07" => data <= "0000000000";
                when x"1C08" => data <= "0000000000";
                when x"1C09" => data <= "0000000000";
                when x"1C0A" => data <= "0000000000";
                when x"1C0B" => data <= "0000000000";
                when x"1C0C" => data <= "0000000000";
                when x"1C0D" => data <= "0000000000";
                when x"1C0E" => data <= "0000000000";
                when x"1C0F" => data <= "0000000000";
                when x"1C10" => data <= "0000000000";
                when x"1C11" => data <= "0111110111";
                when x"1C12" => data <= "0000000000";
                when x"1C13" => data <= "0000000000";
                when x"1C14" => data <= "0000000000";
                when x"1C15" => data <= "0111110111";
                when x"1C16" => data <= "0000000000";
                when x"1C17" => data <= "0000000000";
                when x"1C18" => data <= "0000000000";
                when x"1C19" => data <= "0000000000";
                when x"1C1A" => data <= "0000000000";
                when x"1C1B" => data <= "0000000000";
                when x"1C1C" => data <= "0000000000";
                when x"1C1D" => data <= "0000000000";
                when x"1C1E" => data <= "0000000000";
                when x"1C1F" => data <= "0000000000";
                when x"1C20" => data <= "0000000000";
                when x"1C21" => data <= "0000000000";
                when x"1C22" => data <= "0000000000";
                when x"1C23" => data <= "0000000000";
                when x"1C24" => data <= "0000000000";
                when x"1C25" => data <= "0000000000";
                when x"1C26" => data <= "0000000000";
                when x"1C27" => data <= "0000000000";
                when x"1C28" => data <= "0000000000";
                when x"1C29" => data <= "0000000000";
                when x"1C2A" => data <= "0000000000";
                when x"1C2B" => data <= "0000000000";
                when x"1C2C" => data <= "0000000000";
                when x"1C2D" => data <= "0000000000";
                when x"1C2E" => data <= "0000000000";
                when x"1C2F" => data <= "0000000000";
                when x"1C30" => data <= "0000000000";
                when x"1C31" => data <= "0000000000";
                when x"1C32" => data <= "0000000000";
                when x"1C33" => data <= "0000000000";
                when x"1C34" => data <= "0000000000";
                when x"1C35" => data <= "0000000000";
                when x"1C36" => data <= "0000000000";
                when x"1C37" => data <= "0000000000";
                when x"1C38" => data <= "0000000000";
                when x"1C39" => data <= "0000000000";
                when x"1C3A" => data <= "0000000000";
                when x"1C3B" => data <= "0000000000";
                when x"1C3C" => data <= "0000000000";
                when x"1C3D" => data <= "0000000000";
                when x"1C3E" => data <= "0000000000";
                when x"1C3F" => data <= "0000000000";
                when x"1C40" => data <= "0000000000";
                when x"1C41" => data <= "0000000000";
                when x"1C42" => data <= "0000000000";
                when x"1C43" => data <= "0000000000";
                when x"1C44" => data <= "0000000000";
                when x"1C45" => data <= "0000000000";
                when x"1C46" => data <= "0000000000";
                when x"1C47" => data <= "0000000000";
                when x"1C48" => data <= "0000000000";
                when x"1C49" => data <= "0000000000";
                when x"1C4A" => data <= "0000000000";
                when x"1C4B" => data <= "0000000000";
                when x"1C4C" => data <= "0000000000";
                when x"1C4D" => data <= "0000000000";
                when x"1C4E" => data <= "0000000000";
                when x"1C4F" => data <= "0000000000";
                when x"1C50" => data <= "0000000000";
                when x"1C51" => data <= "0000000000";
                when x"1C52" => data <= "0000000000";
                when x"1C53" => data <= "0000000000";
                when x"1C54" => data <= "0000000000";
                when x"1C55" => data <= "0000000000";
                when x"1C56" => data <= "0000000000";
                when x"1C57" => data <= "0000000000";
                when x"1C58" => data <= "0000000000";
                when x"1C59" => data <= "0000000000";
                when x"1C5A" => data <= "0000000000";
                when x"1C5B" => data <= "0000000000";
                when x"1C5C" => data <= "0000000000";
                when x"1C5D" => data <= "0000000000";
                when x"1C5E" => data <= "0000000000";
                when x"1C5F" => data <= "0000000000";
                when x"1C60" => data <= "0000000000";
                when x"1C61" => data <= "0000000000";
                when x"1C62" => data <= "0000000000";
                when x"1C63" => data <= "0000000000";
                when x"1C64" => data <= "0000000000";
                when x"1C65" => data <= "0000000000";
                when x"1C66" => data <= "0000000000";
                when x"1C67" => data <= "0000000000";
                when x"1C68" => data <= "0000000000";
                when x"1C69" => data <= "0000000000";
                when x"1C6A" => data <= "0000000000";
                when x"1C6B" => data <= "0000000000";
                when x"1C6C" => data <= "0000000000";
                when x"1C6D" => data <= "0000000000";
                when x"1C6E" => data <= "0000000000";
                when x"1C6F" => data <= "0000000000";
                when x"1C70" => data <= "0000000000";
                when x"1C71" => data <= "0000000000";
                when x"1C72" => data <= "0000000000";
                when x"1C73" => data <= "0000000000";
                when x"1C74" => data <= "0000000000";
                when x"1C75" => data <= "0000000000";
                when x"1C76" => data <= "0000000000";
                when x"1C77" => data <= "0011100001";
                when x"1C78" => data <= "0000000000";
                when x"1C79" => data <= "0000000000";
                when x"1C7A" => data <= "0000000000";
                when x"1C7B" => data <= "0000000000";
                when x"1C7C" => data <= "0000000000";
                when x"1C7D" => data <= "0000000000";
                when x"1C7E" => data <= "0000000000";
                when x"1C7F" => data <= "0000000000";
                when x"1C80" => data <= "0000000000";
                when x"1C81" => data <= "0000000000";
                when x"1C82" => data <= "0000000000";
                when x"1C83" => data <= "0000000000";
                when x"1C84" => data <= "0000000000";
                when x"1C85" => data <= "0000000000";
                when x"1C86" => data <= "0000000000";
                when x"1C87" => data <= "0000000000";
                when x"1C88" => data <= "0000000000";
                when x"1C89" => data <= "0000000000";
                when x"1C8A" => data <= "0000000000";
                when x"1C8B" => data <= "0000000000";
                when x"1C8C" => data <= "0000000000";
                when x"1C8D" => data <= "0000000000";
                when x"1C8E" => data <= "0000000000";
                when x"1C8F" => data <= "0000000000";
                when x"1C90" => data <= "0000000000";
                when x"1C91" => data <= "0000000000";
                when x"1C92" => data <= "0000000000";
                when x"1C93" => data <= "0000000000";
                when x"1C94" => data <= "0000000000";
                when x"1C95" => data <= "0000000000";
                when x"1C96" => data <= "0000000000";
                when x"1C97" => data <= "0000000000";
                when x"1C98" => data <= "0000000000";
                when x"1C99" => data <= "0000000000";
                when x"1C9A" => data <= "0000000000";
                when x"1C9B" => data <= "0000000000";
                when x"1C9C" => data <= "0000000000";
                when x"1C9D" => data <= "0000000000";
                when x"1C9E" => data <= "0000000000";
                when x"1C9F" => data <= "0000000000";
                when x"1CA0" => data <= "0000000000";
                when x"1CA1" => data <= "0000000000";
                when x"1CA2" => data <= "0000000000";
                when x"1CA3" => data <= "0000000000";
                when x"1CA4" => data <= "0000000000";
                when x"1CA5" => data <= "0000000000";
                when x"1CA6" => data <= "0000000000";
                when x"1CA7" => data <= "0000000000";
                when x"1CA8" => data <= "0000000000";
                when x"1CA9" => data <= "0000000000";
                when x"1CAA" => data <= "0000000000";
                when x"1CAB" => data <= "0000000000";
                when x"1CAC" => data <= "0000000000";
                when x"1CAD" => data <= "0000000000";
                when x"1CAE" => data <= "0000000000";
                when x"1CAF" => data <= "0000000000";
                when x"1CB0" => data <= "0000000000";
                when x"1CB1" => data <= "0000000000";
                when x"1CB2" => data <= "0000000000";
                when x"1CB3" => data <= "0000000000";
                when x"1CB4" => data <= "0000000000";
                when x"1CB5" => data <= "0000000000";
                when x"1CB6" => data <= "0000000000";
                when x"1CB7" => data <= "0000000000";
                when x"1CB8" => data <= "0000000000";
                when x"1CB9" => data <= "0000000000";
                when x"1CBA" => data <= "0000000000";
                when x"1CBB" => data <= "0000000000";
                when x"1CBC" => data <= "0000000000";
                when x"1CBD" => data <= "0000000000";
                when x"1CBE" => data <= "0000000000";
                when x"1CBF" => data <= "0000000000";
                when x"1CC0" => data <= "0000000000";
                when x"1CC1" => data <= "0000000000";
                when x"1CC2" => data <= "0000000000";
                when x"1CC3" => data <= "0000000000";
                when x"1CC4" => data <= "0000000000";
                when x"1CC5" => data <= "0000000000";
                when x"1CC6" => data <= "0000000000";
                when x"1CC7" => data <= "0000000000";
                when x"1CC8" => data <= "0000000000";
                when x"1CC9" => data <= "0000000000";
                when x"1CCA" => data <= "0000000000";
                when x"1CCB" => data <= "0000000000";
                when x"1CCC" => data <= "0000000000";
                when x"1CCD" => data <= "0000000000";
                when x"1CCE" => data <= "0000000000";
                when x"1CCF" => data <= "0000000000";
                when x"1CD0" => data <= "0000000000";
                when x"1CD1" => data <= "0000000000";
                when x"1CD2" => data <= "0000000000";
                when x"1CD3" => data <= "0000000000";
                when x"1CD4" => data <= "0000000000";
                when x"1CD5" => data <= "0000000000";
                when x"1CD6" => data <= "0000000000";
                when x"1CD7" => data <= "0000000000";
                when x"1CD8" => data <= "0000000000";
                when x"1CD9" => data <= "0000000000";
                when x"1CDA" => data <= "0000000000";
                when x"1CDB" => data <= "0000000000";
                when x"1CDC" => data <= "0000000000";
                when x"1CDD" => data <= "0000000000";
                when x"1CDE" => data <= "0000000000";
                when x"1CDF" => data <= "0000000000";
                when x"1CE0" => data <= "0000000000";
                when x"1CE1" => data <= "0000000000";
                when x"1CE2" => data <= "0000000000";
                when x"1CE3" => data <= "0000000000";
                when x"1CE4" => data <= "0000000000";
                when x"1CE5" => data <= "0000000000";
                when x"1CE6" => data <= "0000000000";
                when x"1CE7" => data <= "0000000000";
                when x"1CE8" => data <= "0000000000";
                when x"1CE9" => data <= "0000000000";
                when x"1CEA" => data <= "0000000000";
                when x"1CEB" => data <= "0000000000";
                when x"1CEC" => data <= "0000000000";
                when x"1CED" => data <= "0000000000";
                when x"1CEE" => data <= "0000000000";
                when x"1CEF" => data <= "0000000000";
                when x"1CF0" => data <= "0000000000";
                when x"1CF1" => data <= "0000000000";
                when x"1CF2" => data <= "0000000000";
                when x"1CF3" => data <= "0000000000";
                when x"1CF4" => data <= "0000000000";
                when x"1CF5" => data <= "0000000000";
                when x"1CF6" => data <= "0000000000";
                when x"1CF7" => data <= "0000000000";
                when x"1CF8" => data <= "0000000000";
                when x"1CF9" => data <= "0000000000";
                when x"1CFA" => data <= "0000000000";
                when x"1CFB" => data <= "0000000000";
                when x"1CFC" => data <= "0000000000";
                when x"1CFD" => data <= "0000000000";
                when x"1CFE" => data <= "0000000000";
                when x"1CFF" => data <= "0000000000";
                when x"1D00" => data <= "0000000000";
                when x"1D01" => data <= "0000000000";
                when x"1D02" => data <= "0000000000";
                when x"1D03" => data <= "0000000000";
                when x"1D04" => data <= "0000000000";
                when x"1D05" => data <= "0000000000";
                when x"1D06" => data <= "0000000000";
                when x"1D07" => data <= "0000000000";
                when x"1D08" => data <= "0000000000";
                when x"1D09" => data <= "0000000000";
                when x"1D0A" => data <= "0000000000";
                when x"1D0B" => data <= "0000000000";
                when x"1D0C" => data <= "0000000000";
                when x"1D0D" => data <= "0000000000";
                when x"1D0E" => data <= "0000000000";
                when x"1D0F" => data <= "0000000000";
                when x"1D10" => data <= "1000101100";
                when x"1D11" => data <= "0000000000";
                when x"1D12" => data <= "0000000000";
                when x"1D13" => data <= "0000000000";
                when x"1D14" => data <= "0000000000";
                when x"1D15" => data <= "0000000000";
                when x"1D16" => data <= "0000000000";
                when x"1D17" => data <= "0000000000";
                when x"1D18" => data <= "0000000000";
                when x"1D19" => data <= "0000000000";
                when x"1D1A" => data <= "0000000000";
                when x"1D1B" => data <= "0000000000";
                when x"1D1C" => data <= "0000000000";
                when x"1D1D" => data <= "0000000000";
                when x"1D1E" => data <= "0000000000";
                when x"1D1F" => data <= "0000000000";
                when x"1D20" => data <= "0000000000";
                when x"1D21" => data <= "0000000000";
                when x"1D22" => data <= "0000000000";
                when x"1D23" => data <= "0000000000";
                when x"1D24" => data <= "0000000000";
                when x"1D25" => data <= "0000000000";
                when x"1D26" => data <= "0000000000";
                when x"1D27" => data <= "0000000000";
                when x"1D28" => data <= "0000000000";
                when x"1D29" => data <= "0000000000";
                when x"1D2A" => data <= "0000000000";
                when x"1D2B" => data <= "0000000000";
                when x"1D2C" => data <= "0000000000";
                when x"1D2D" => data <= "0000000000";
                when x"1D2E" => data <= "0000000000";
                when x"1D2F" => data <= "0000000000";
                when x"1D30" => data <= "0000000000";
                when x"1D31" => data <= "0000000000";
                when x"1D32" => data <= "0000000000";
                when x"1D33" => data <= "0000000000";
                when x"1D34" => data <= "0000000000";
                when x"1D35" => data <= "0000000000";
                when x"1D36" => data <= "1111011011";
                when x"1D37" => data <= "0000000000";
                when x"1D38" => data <= "0000000000";
                when x"1D39" => data <= "0000000000";
                when x"1D3A" => data <= "0000000000";
                when x"1D3B" => data <= "0000000000";
                when x"1D3C" => data <= "0000000000";
                when x"1D3D" => data <= "0000000000";
                when x"1D3E" => data <= "0000000000";
                when x"1D3F" => data <= "0000000000";
                when x"1D40" => data <= "0000000000";
                when x"1D41" => data <= "0000000000";
                when x"1D42" => data <= "0000000000";
                when x"1D43" => data <= "0000000000";
                when x"1D44" => data <= "0000000000";
                when x"1D45" => data <= "0000000000";
                when x"1D46" => data <= "0000000000";
                when x"1D47" => data <= "0000000000";
                when x"1D48" => data <= "0000000000";
                when x"1D49" => data <= "0000000000";
                when x"1D4A" => data <= "0000000000";
                when x"1D4B" => data <= "0000000000";
                when x"1D4C" => data <= "0000000000";
                when x"1D4D" => data <= "0000000000";
                when x"1D4E" => data <= "0000000000";
                when x"1D4F" => data <= "0000000000";
                when x"1D50" => data <= "0000000000";
                when x"1D51" => data <= "0000000000";
                when x"1D52" => data <= "0000000000";
                when x"1D53" => data <= "0000000000";
                when x"1D54" => data <= "0000000000";
                when x"1D55" => data <= "0000000000";
                when x"1D56" => data <= "1111011011";
                when x"1D57" => data <= "0000000000";
                when x"1D58" => data <= "0000000000";
                when x"1D59" => data <= "0000000000";
                when x"1D5A" => data <= "0000000000";
                when x"1D5B" => data <= "0000000000";
                when x"1D5C" => data <= "0000000000";
                when x"1D5D" => data <= "0000000000";
                when x"1D5E" => data <= "0000000000";
                when x"1D5F" => data <= "0000000000";
                when x"1D60" => data <= "0000000000";
                when x"1D61" => data <= "0000000000";
                when x"1D62" => data <= "0000000000";
                when x"1D63" => data <= "0000000000";
                when x"1D64" => data <= "0000000000";
                when x"1D65" => data <= "0000000000";
                when x"1D66" => data <= "0000000000";
                when x"1D67" => data <= "0000000000";
                when x"1D68" => data <= "0000000000";
                when x"1D69" => data <= "1111011011";
                when x"1D6A" => data <= "0000000000";
                when x"1D6B" => data <= "0000000000";
                when x"1D6C" => data <= "0000000000";
                when x"1D6D" => data <= "0000000000";
                when x"1D6E" => data <= "0000000000";
                when x"1D6F" => data <= "0000000000";
                when x"1D70" => data <= "0000000000";
                when x"1D71" => data <= "0000000000";
                when x"1D72" => data <= "0000000000";
                when x"1D73" => data <= "0000000000";
                when x"1D74" => data <= "0000000000";
                when x"1D75" => data <= "0000000000";
                when x"1D76" => data <= "0000000000";
                when x"1D77" => data <= "0000000000";
                when x"1D78" => data <= "0000000000";
                when x"1D79" => data <= "0000000000";
                when x"1D7A" => data <= "0000000000";
                when x"1D7B" => data <= "0000000000";
                when x"1D7C" => data <= "0000000000";
                when x"1D7D" => data <= "0100100011";
                when x"1D7E" => data <= "0000000000";
                when x"1D7F" => data <= "0000000000";
                when x"1D80" => data <= "0000000000";
                when x"1D81" => data <= "0000000000";
                when x"1D82" => data <= "0000000000";
                when x"1D83" => data <= "0000000000";
                when x"1D84" => data <= "0000000000";
                when x"1D85" => data <= "0000000000";
                when x"1D86" => data <= "0000000000";
                when x"1D87" => data <= "0000000000";
                when x"1D88" => data <= "0000000000";
                when x"1D89" => data <= "0000000000";
                when x"1D8A" => data <= "0000000000";
                when x"1D8B" => data <= "0000000000";
                when x"1D8C" => data <= "0000000000";
                when x"1D8D" => data <= "0000000000";
                when x"1D8E" => data <= "0000000000";
                when x"1D8F" => data <= "0000000000";
                when x"1D90" => data <= "0000000000";
                when x"1D91" => data <= "0000000000";
                when x"1D92" => data <= "0000000000";
                when x"1D93" => data <= "0000000000";
                when x"1D94" => data <= "0000000000";
                when x"1D95" => data <= "0000000000";
                when x"1D96" => data <= "0000000000";
                when x"1D97" => data <= "0000000000";
                when x"1D98" => data <= "0000000000";
                when x"1D99" => data <= "0000000000";
                when x"1D9A" => data <= "0000000000";
                when x"1D9B" => data <= "0000000000";
                when x"1D9C" => data <= "0000000000";
                when x"1D9D" => data <= "0000000000";
                when x"1D9E" => data <= "0000000000";
                when x"1D9F" => data <= "0000000000";
                when x"1DA0" => data <= "0000000000";
                when x"1DA1" => data <= "0000000000";
                when x"1DA2" => data <= "0000000000";
                when x"1DA3" => data <= "0000000000";
                when x"1DA4" => data <= "0000000000";
                when x"1DA5" => data <= "0000000000";
                when x"1DA6" => data <= "0000000000";
                when x"1DA7" => data <= "0000000000";
                when x"1DA8" => data <= "0000000000";
                when x"1DA9" => data <= "0000000000";
                when x"1DAA" => data <= "0000000000";
                when x"1DAB" => data <= "0000000000";
                when x"1DAC" => data <= "0000000000";
                when x"1DAD" => data <= "0000000000";
                when x"1DAE" => data <= "0000000000";
                when x"1DAF" => data <= "0000000000";
                when x"1DB0" => data <= "0000000000";
                when x"1DB1" => data <= "0000000000";
                when x"1DB2" => data <= "0000000000";
                when x"1DB3" => data <= "0000000000";
                when x"1DB4" => data <= "0000000000";
                when x"1DB5" => data <= "0000000000";
                when x"1DB6" => data <= "0000000000";
                when x"1DB7" => data <= "0000000000";
                when x"1DB8" => data <= "0000000000";
                when x"1DB9" => data <= "0000000000";
                when x"1DBA" => data <= "0000000000";
                when x"1DBB" => data <= "0000000000";
                when x"1DBC" => data <= "0000000000";
                when x"1DBD" => data <= "0000000000";
                when x"1DBE" => data <= "0000000000";
                when x"1DBF" => data <= "0000000000";
                when x"1DC0" => data <= "0000000000";
                when x"1DC1" => data <= "0000000000";
                when x"1DC2" => data <= "0000000000";
                when x"1DC3" => data <= "0000000000";
                when x"1DC4" => data <= "0000000000";
                when x"1DC5" => data <= "0000000000";
                when x"1DC6" => data <= "0000000000";
                when x"1DC7" => data <= "0000000000";
                when x"1DC8" => data <= "0000000000";
                when x"1DC9" => data <= "0000000000";
                when x"1DCA" => data <= "0000000000";
                when x"1DCB" => data <= "0000000000";
                when x"1DCC" => data <= "0000000000";
                when x"1DCD" => data <= "0000000000";
                when x"1DCE" => data <= "1011001101";
                when x"1DCF" => data <= "0000000000";
                when x"1DD0" => data <= "0000000000";
                when x"1DD1" => data <= "0000000000";
                when x"1DD2" => data <= "0000000000";
                when x"1DD3" => data <= "0000000000";
                when x"1DD4" => data <= "0000000000";
                when x"1DD5" => data <= "0000000000";
                when x"1DD6" => data <= "0000000000";
                when x"1DD7" => data <= "0000000000";
                when x"1DD8" => data <= "0000000000";
                when x"1DD9" => data <= "0000000000";
                when x"1DDA" => data <= "0000000000";
                when x"1DDB" => data <= "0000000000";
                when x"1DDC" => data <= "0000000000";
                when x"1DDD" => data <= "0000000000";
                when x"1DDE" => data <= "0000000000";
                when x"1DDF" => data <= "0000000000";
                when x"1DE0" => data <= "0000000000";
                when x"1DE1" => data <= "0000000000";
                when x"1DE2" => data <= "0000000000";
                when x"1DE3" => data <= "0000000000";
                when x"1DE4" => data <= "0000000000";
                when x"1DE5" => data <= "0000000000";
                when x"1DE6" => data <= "0000000000";
                when x"1DE7" => data <= "0000000000";
                when x"1DE8" => data <= "0000000000";
                when x"1DE9" => data <= "0000000000";
                when x"1DEA" => data <= "0000000000";
                when x"1DEB" => data <= "0000000000";
                when x"1DEC" => data <= "0000000000";
                when x"1DED" => data <= "0000000000";
                when x"1DEE" => data <= "0000000000";
                when x"1DEF" => data <= "0000000000";
                when x"1DF0" => data <= "0000000000";
                when x"1DF1" => data <= "0000000000";
                when x"1DF2" => data <= "0000000000";
                when x"1DF3" => data <= "0000000000";
                when x"1DF4" => data <= "0000000000";
                when x"1DF5" => data <= "0000000000";
                when x"1DF6" => data <= "0000000000";
                when x"1DF7" => data <= "0000000000";
                when x"1DF8" => data <= "0000000000";
                when x"1DF9" => data <= "0000000000";
                when x"1DFA" => data <= "0000000000";
                when x"1DFB" => data <= "0000000000";
                when x"1DFC" => data <= "0000000000";
                when x"1DFD" => data <= "0000000000";
                when x"1DFE" => data <= "0000000000";
                when x"1DFF" => data <= "0000000000";
                when x"1E00" => data <= "0000000000";
                when x"1E01" => data <= "0000000000";
                when x"1E02" => data <= "0000000000";
                when x"1E03" => data <= "0000000000";
                when x"1E04" => data <= "0000000000";
                when x"1E05" => data <= "0000000000";
                when x"1E06" => data <= "0000000000";
                when x"1E07" => data <= "0000000000";
                when x"1E08" => data <= "0000000000";
                when x"1E09" => data <= "0000000000";
                when x"1E0A" => data <= "0000000000";
                when x"1E0B" => data <= "0000000000";
                when x"1E0C" => data <= "0000000000";
                when x"1E0D" => data <= "0000000000";
                when x"1E0E" => data <= "0000000000";
                when x"1E0F" => data <= "0000000000";
                when x"1E10" => data <= "0000000000";
                when x"1E11" => data <= "0000000000";
                when x"1E12" => data <= "0111110111";
                when x"1E13" => data <= "0000000000";
                when x"1E14" => data <= "0000000000";
                when x"1E15" => data <= "0000000000";
                when x"1E16" => data <= "0000000000";
                when x"1E17" => data <= "0000000000";
                when x"1E18" => data <= "0000000000";
                when x"1E19" => data <= "0000000000";
                when x"1E1A" => data <= "0000000000";
                when x"1E1B" => data <= "0000000000";
                when x"1E1C" => data <= "0000000000";
                when x"1E1D" => data <= "0000000000";
                when x"1E1E" => data <= "0000000000";
                when x"1E1F" => data <= "0000000000";
                when x"1E20" => data <= "0000000000";
                when x"1E21" => data <= "0000000000";
                when x"1E22" => data <= "0000000000";
                when x"1E23" => data <= "0000000000";
                when x"1E24" => data <= "0000000000";
                when x"1E25" => data <= "0000000000";
                when x"1E26" => data <= "0000000000";
                when x"1E27" => data <= "0000000000";
                when x"1E28" => data <= "0000000000";
                when x"1E29" => data <= "0000000000";
                when x"1E2A" => data <= "0000000000";
                when x"1E2B" => data <= "0000000000";
                when x"1E2C" => data <= "0000000000";
                when x"1E2D" => data <= "0000000000";
                when x"1E2E" => data <= "0000000000";
                when x"1E2F" => data <= "0000000000";
                when x"1E30" => data <= "0000000000";
                when x"1E31" => data <= "0000000000";
                when x"1E32" => data <= "0000000000";
                when x"1E33" => data <= "0000000000";
                when x"1E34" => data <= "0000000000";
                when x"1E35" => data <= "0000000000";
                when x"1E36" => data <= "0000000000";
                when x"1E37" => data <= "0000000000";
                when x"1E38" => data <= "0000000000";
                when x"1E39" => data <= "0000000000";
                when x"1E3A" => data <= "0000000000";
                when x"1E3B" => data <= "0000000000";
                when x"1E3C" => data <= "0000000000";
                when x"1E3D" => data <= "0000000000";
                when x"1E3E" => data <= "0000000000";
                when x"1E3F" => data <= "0000000000";
                when x"1E40" => data <= "0000000000";
                when x"1E41" => data <= "0000000000";
                when x"1E42" => data <= "0000000000";
                when x"1E43" => data <= "0000000000";
                when x"1E44" => data <= "0000000000";
                when x"1E45" => data <= "0000000000";
                when x"1E46" => data <= "0000000000";
                when x"1E47" => data <= "0000000000";
                when x"1E48" => data <= "0000000000";
                when x"1E49" => data <= "0000000000";
                when x"1E4A" => data <= "1101010000";
                when x"1E4B" => data <= "0000000000";
                when x"1E4C" => data <= "0000000000";
                when x"1E4D" => data <= "0000000000";
                when x"1E4E" => data <= "0000000000";
                when x"1E4F" => data <= "0000000000";
                when x"1E50" => data <= "0000000000";
                when x"1E51" => data <= "0000000000";
                when x"1E52" => data <= "0000000000";
                when x"1E53" => data <= "0000000000";
                when x"1E54" => data <= "0000000000";
                when x"1E55" => data <= "0000000000";
                when x"1E56" => data <= "0000000000";
                when x"1E57" => data <= "0000000000";
                when x"1E58" => data <= "0000000000";
                when x"1E59" => data <= "0000000000";
                when x"1E5A" => data <= "0000000000";
                when x"1E5B" => data <= "0000000000";
                when x"1E5C" => data <= "0000000000";
                when x"1E5D" => data <= "0000000000";
                when x"1E5E" => data <= "0000000000";
                when x"1E5F" => data <= "0000000000";
                when x"1E60" => data <= "0000000000";
                when x"1E61" => data <= "0000000000";
                when x"1E62" => data <= "0000000000";
                when x"1E63" => data <= "0000000000";
                when x"1E64" => data <= "0000000000";
                when x"1E65" => data <= "0000000000";
                when x"1E66" => data <= "0000000000";
                when x"1E67" => data <= "0000000000";
                when x"1E68" => data <= "0000000000";
                when x"1E69" => data <= "0000000000";
                when x"1E6A" => data <= "0000000000";
                when x"1E6B" => data <= "0000000000";
                when x"1E6C" => data <= "0000000000";
                when x"1E6D" => data <= "0000000000";
                when x"1E6E" => data <= "0000000000";
                when x"1E6F" => data <= "0000000000";
                when x"1E70" => data <= "0000000000";
                when x"1E71" => data <= "0000000000";
                when x"1E72" => data <= "0000000000";
                when x"1E73" => data <= "0000000000";
                when x"1E74" => data <= "0000000000";
                when x"1E75" => data <= "0000000000";
                when x"1E76" => data <= "0000000000";
                when x"1E77" => data <= "0000000000";
                when x"1E78" => data <= "0000000000";
                when x"1E79" => data <= "0000000000";
                when x"1E7A" => data <= "0000000000";
                when x"1E7B" => data <= "0000000000";
                when x"1E7C" => data <= "0000000000";
                when x"1E7D" => data <= "0000000000";
                when x"1E7E" => data <= "0000000000";
                when x"1E7F" => data <= "0000000000";
                when x"1E80" => data <= "0000000000";
                when x"1E81" => data <= "0000000000";
                when x"1E82" => data <= "0000000000";
                when x"1E83" => data <= "0000000000";
                when x"1E84" => data <= "0000000000";
                when x"1E85" => data <= "0000000000";
                when x"1E86" => data <= "0000000000";
                when x"1E87" => data <= "0000000000";
                when x"1E88" => data <= "0000000000";
                when x"1E89" => data <= "0000000000";
                when x"1E8A" => data <= "0000000000";
                when x"1E8B" => data <= "0000000000";
                when x"1E8C" => data <= "0000000000";
                when x"1E8D" => data <= "0000000000";
                when x"1E8E" => data <= "0000000000";
                when x"1E8F" => data <= "0000000000";
                when x"1E90" => data <= "0000000000";
                when x"1E91" => data <= "0000000000";
                when x"1E92" => data <= "0000000000";
                when x"1E93" => data <= "0000000000";
                when x"1E94" => data <= "0000000000";
                when x"1E95" => data <= "0000000000";
                when x"1E96" => data <= "0000000000";
                when x"1E97" => data <= "0000000000";
                when x"1E98" => data <= "0000000000";
                when x"1E99" => data <= "0000000000";
                when x"1E9A" => data <= "0000000000";
                when x"1E9B" => data <= "0000000000";
                when x"1E9C" => data <= "0000000000";
                when x"1E9D" => data <= "0000000000";
                when x"1E9E" => data <= "0000000000";
                when x"1E9F" => data <= "0000000000";
                when x"1EA0" => data <= "0000000000";
                when x"1EA1" => data <= "0000000000";
                when x"1EA2" => data <= "0000000000";
                when x"1EA3" => data <= "0000000000";
                when x"1EA4" => data <= "0000000000";
                when x"1EA5" => data <= "0000000000";
                when x"1EA6" => data <= "0000000000";
                when x"1EA7" => data <= "0000000000";
                when x"1EA8" => data <= "0000000000";
                when x"1EA9" => data <= "0000000000";
                when x"1EAA" => data <= "0000000000";
                when x"1EAB" => data <= "0000000000";
                when x"1EAC" => data <= "0000000000";
                when x"1EAD" => data <= "0111110111";
                when x"1EAE" => data <= "0000000000";
                when x"1EAF" => data <= "0000000000";
                when x"1EB0" => data <= "0000000000";
                when x"1EB1" => data <= "0000000000";
                when x"1EB2" => data <= "0000000000";
                when x"1EB3" => data <= "0000000000";
                when x"1EB4" => data <= "0000000000";
                when x"1EB5" => data <= "0000000000";
                when x"1EB6" => data <= "0000000000";
                when x"1EB7" => data <= "0000000000";
                when x"1EB8" => data <= "0000000000";
                when x"1EB9" => data <= "0000000000";
                when x"1EBA" => data <= "0000000000";
                when x"1EBB" => data <= "0000000000";
                when x"1EBC" => data <= "0000000000";
                when x"1EBD" => data <= "0000000000";
                when x"1EBE" => data <= "0000000000";
                when x"1EBF" => data <= "0000000000";
                when x"1EC0" => data <= "0000000000";
                when x"1EC1" => data <= "0000000000";
                when x"1EC2" => data <= "0000000000";
                when x"1EC3" => data <= "0000000000";
                when x"1EC4" => data <= "0000000000";
                when x"1EC5" => data <= "0000000000";
                when x"1EC6" => data <= "0000000000";
                when x"1EC7" => data <= "0000000000";
                when x"1EC8" => data <= "0000000000";
                when x"1EC9" => data <= "0000000000";
                when x"1ECA" => data <= "0000000000";
                when x"1ECB" => data <= "0000000000";
                when x"1ECC" => data <= "0000000000";
                when x"1ECD" => data <= "0000000000";
                when x"1ECE" => data <= "0000000000";
                when x"1ECF" => data <= "0000000000";
                when x"1ED0" => data <= "0000000000";
                when x"1ED1" => data <= "0000000000";
                when x"1ED2" => data <= "0000000000";
                when x"1ED3" => data <= "0000000000";
                when x"1ED4" => data <= "0000000000";
                when x"1ED5" => data <= "0000000000";
                when x"1ED6" => data <= "0000000000";
                when x"1ED7" => data <= "0000000000";
                when x"1ED8" => data <= "0000000000";
                when x"1ED9" => data <= "0000000000";
                when x"1EDA" => data <= "0000000000";
                when x"1EDB" => data <= "0000000000";
                when x"1EDC" => data <= "0000000000";
                when x"1EDD" => data <= "0000000000";
                when x"1EDE" => data <= "0000000000";
                when x"1EDF" => data <= "0000000000";
                when x"1EE0" => data <= "0000000000";
                when x"1EE1" => data <= "0000000000";
                when x"1EE2" => data <= "0000000000";
                when x"1EE3" => data <= "0000000000";
                when x"1EE4" => data <= "0000000000";
                when x"1EE5" => data <= "0000000000";
                when x"1EE6" => data <= "0000000000";
                when x"1EE7" => data <= "0000000000";
                when x"1EE8" => data <= "0000000000";
                when x"1EE9" => data <= "0000000000";
                when x"1EEA" => data <= "0000000000";
                when x"1EEB" => data <= "0000000000";
                when x"1EEC" => data <= "0000000000";
                when x"1EED" => data <= "0000000000";
                when x"1EEE" => data <= "0000000000";
                when x"1EEF" => data <= "0000000000";
                when x"1EF0" => data <= "0000000000";
                when x"1EF1" => data <= "0000000000";
                when x"1EF2" => data <= "0000000000";
                when x"1EF3" => data <= "0000000000";
                when x"1EF4" => data <= "0000000000";
                when x"1EF5" => data <= "0000000000";
                when x"1EF6" => data <= "0000000000";
                when x"1EF7" => data <= "0000000000";
                when x"1EF8" => data <= "0000000000";
                when x"1EF9" => data <= "0000000000";
                when x"1EFA" => data <= "0000000000";
                when x"1EFB" => data <= "0000000000";
                when x"1EFC" => data <= "0000000000";
                when x"1EFD" => data <= "0000000000";
                when x"1EFE" => data <= "0000000000";
                when x"1EFF" => data <= "0000000000";
                when x"1F00" => data <= "0000000000";
                when x"1F01" => data <= "0000000000";
                when x"1F02" => data <= "0000000000";
                when x"1F03" => data <= "0000000000";
                when x"1F04" => data <= "0000000000";
                when x"1F05" => data <= "0000000000";
                when x"1F06" => data <= "0000000000";
                when x"1F07" => data <= "0000000000";
                when x"1F08" => data <= "0000000000";
                when x"1F09" => data <= "0000000000";
                when x"1F0A" => data <= "0000000000";
                when x"1F0B" => data <= "0000000000";
                when x"1F0C" => data <= "0000000000";
                when x"1F0D" => data <= "0000000000";
                when x"1F0E" => data <= "0000000000";
                when x"1F0F" => data <= "0000000000";
                when x"1F10" => data <= "0000000000";
                when x"1F11" => data <= "0000000000";
                when x"1F12" => data <= "0000000000";
                when x"1F13" => data <= "0000000000";
                when x"1F14" => data <= "0000000000";
                when x"1F15" => data <= "0000000000";
                when x"1F16" => data <= "0000000000";
                when x"1F17" => data <= "0000000000";
                when x"1F18" => data <= "0000000000";
                when x"1F19" => data <= "0000000000";
                when x"1F1A" => data <= "0000000000";
                when x"1F1B" => data <= "0000000000";
                when x"1F1C" => data <= "0000000000";
                when x"1F1D" => data <= "0000000000";
                when x"1F1E" => data <= "0000000000";
                when x"1F1F" => data <= "0000000000";
                when x"1F20" => data <= "0000000000";
                when x"1F21" => data <= "0000000000";
                when x"1F22" => data <= "0000000000";
                when x"1F23" => data <= "0000000000";
                when x"1F24" => data <= "0000000000";
                when x"1F25" => data <= "0000000000";
                when x"1F26" => data <= "0000000000";
                when x"1F27" => data <= "0000000000";
                when x"1F28" => data <= "0000000000";
                when x"1F29" => data <= "0000000000";
                when x"1F2A" => data <= "0000000000";
                when x"1F2B" => data <= "0000000000";
                when x"1F2C" => data <= "0000000000";
                when x"1F2D" => data <= "0000000000";
                when x"1F2E" => data <= "0000000000";
                when x"1F2F" => data <= "0000000000";
                when x"1F30" => data <= "0000000000";
                when x"1F31" => data <= "0000000000";
                when x"1F32" => data <= "0000000000";
                when x"1F33" => data <= "0000000000";
                when x"1F34" => data <= "0000000000";
                when x"1F35" => data <= "0000000000";
                when x"1F36" => data <= "0000000000";
                when x"1F37" => data <= "0000000000";
                when x"1F38" => data <= "0000000000";
                when x"1F39" => data <= "0000000000";
                when x"1F3A" => data <= "0000000000";
                when x"1F3B" => data <= "0000000000";
                when x"1F3C" => data <= "0000000000";
                when x"1F3D" => data <= "0000000000";
                when x"1F3E" => data <= "0000000000";
                when x"1F3F" => data <= "0000000000";
                when x"1F40" => data <= "0000000000";
                when x"1F41" => data <= "0000000000";
                when x"1F42" => data <= "0000000000";
                when x"1F43" => data <= "0000000000";
                when x"1F44" => data <= "0000000000";
                when x"1F45" => data <= "0000000000";
                when x"1F46" => data <= "0000000000";
                when x"1F47" => data <= "0000000000";
                when x"1F48" => data <= "0000000000";
                when x"1F49" => data <= "0000000000";
                when x"1F4A" => data <= "0000000000";
                when x"1F4B" => data <= "0000000000";
                when x"1F4C" => data <= "0000000000";
                when x"1F4D" => data <= "0000000000";
                when x"1F4E" => data <= "0000000000";
                when x"1F4F" => data <= "0000000000";
                when x"1F50" => data <= "0000000000";
                when x"1F51" => data <= "0000000000";
                when x"1F52" => data <= "0000000000";
                when x"1F53" => data <= "0000000000";
                when x"1F54" => data <= "0000000000";
                when x"1F55" => data <= "0000000000";
                when x"1F56" => data <= "0000000000";
                when x"1F57" => data <= "0000000000";
                when x"1F58" => data <= "0000000000";
                when x"1F59" => data <= "0000000000";
                when x"1F5A" => data <= "0000000000";
                when x"1F5B" => data <= "0000000000";
                when x"1F5C" => data <= "0000000000";
                when x"1F5D" => data <= "0000000000";
                when x"1F5E" => data <= "0000000000";
                when x"1F5F" => data <= "0000000000";
                when x"1F60" => data <= "0000000000";
                when x"1F61" => data <= "0000000000";
                when x"1F62" => data <= "0000000000";
                when x"1F63" => data <= "0000000000";
                when x"1F64" => data <= "0000000000";
                when x"1F65" => data <= "0000000000";
                when x"1F66" => data <= "0000000000";
                when x"1F67" => data <= "0000000000";
                when x"1F68" => data <= "0111000010";
                when x"1F69" => data <= "0000000000";
                when x"1F6A" => data <= "0000000000";
                when x"1F6B" => data <= "0000000000";
                when x"1F6C" => data <= "0000000000";
                when x"1F6D" => data <= "0000000000";
                when x"1F6E" => data <= "0000000000";
                when x"1F6F" => data <= "0000000000";
                when x"1F70" => data <= "0000000000";
                when x"1F71" => data <= "0000000000";
                when x"1F72" => data <= "0000000000";
                when x"1F73" => data <= "0000000000";
                when x"1F74" => data <= "0000000000";
                when x"1F75" => data <= "0000000000";
                when x"1F76" => data <= "0000000000";
                when x"1F77" => data <= "0000000000";
                when x"1F78" => data <= "0000000000";
                when x"1F79" => data <= "0000000000";
                when x"1F7A" => data <= "0000000000";
                when x"1F7B" => data <= "0000000000";
                when x"1F7C" => data <= "0000000000";
                when x"1F7D" => data <= "0000000000";
                when x"1F7E" => data <= "0000000000";
                when x"1F7F" => data <= "0000000000";
                when x"1F80" => data <= "0000000000";
                when x"1F81" => data <= "0000000000";
                when x"1F82" => data <= "0000000000";
                when x"1F83" => data <= "0000000000";
                when x"1F84" => data <= "0000000000";
                when x"1F85" => data <= "0000000000";
                when x"1F86" => data <= "0000000000";
                when x"1F87" => data <= "0000000000";
                when x"1F88" => data <= "0000000000";
                when x"1F89" => data <= "0000000000";
                when x"1F8A" => data <= "0000000000";
                when x"1F8B" => data <= "0000000000";
                when x"1F8C" => data <= "0000000000";
                when x"1F8D" => data <= "0000000000";
                when x"1F8E" => data <= "0000000000";
                when x"1F8F" => data <= "0000000000";
                when x"1F90" => data <= "0111110111";
                when x"1F91" => data <= "0000000000";
                when x"1F92" => data <= "0000000000";
                when x"1F93" => data <= "0000000000";
                when x"1F94" => data <= "0000000000";
                when x"1F95" => data <= "0000000000";
                when x"1F96" => data <= "0000000000";
                when x"1F97" => data <= "0000000000";
                when x"1F98" => data <= "0000000000";
                when x"1F99" => data <= "0000000000";
                when x"1F9A" => data <= "0000000000";
                when x"1F9B" => data <= "0000000000";
                when x"1F9C" => data <= "0000000000";
                when x"1F9D" => data <= "0000000000";
                when x"1F9E" => data <= "0000000000";
                when x"1F9F" => data <= "0000000000";
                when x"1FA0" => data <= "0000000000";
                when x"1FA1" => data <= "0000000000";
                when x"1FA2" => data <= "0000000000";
                when x"1FA3" => data <= "0000000000";
                when x"1FA4" => data <= "0000000000";
                when x"1FA5" => data <= "0000000000";
                when x"1FA6" => data <= "0000000000";
                when x"1FA7" => data <= "0000000000";
                when x"1FA8" => data <= "0000000000";
                when x"1FA9" => data <= "0000000000";
                when x"1FAA" => data <= "0000000000";
                when x"1FAB" => data <= "0000000000";
                when x"1FAC" => data <= "0000000000";
                when x"1FAD" => data <= "0000000000";
                when x"1FAE" => data <= "0000000000";
                when x"1FAF" => data <= "0000000000";
                when x"1FB0" => data <= "0000000000";
                when x"1FB1" => data <= "0000000000";
                when x"1FB2" => data <= "0000000000";
                when x"1FB3" => data <= "0000000000";
                when x"1FB4" => data <= "0000000000";
                when x"1FB5" => data <= "0000000000";
                when x"1FB6" => data <= "0000000000";
                when x"1FB7" => data <= "0000000000";
                when x"1FB8" => data <= "0000000000";
                when x"1FB9" => data <= "0000000000";
                when x"1FBA" => data <= "0000000000";
                when x"1FBB" => data <= "0000000000";
                when x"1FBC" => data <= "0000000000";
                when x"1FBD" => data <= "0000000000";
                when x"1FBE" => data <= "0000000000";
                when x"1FBF" => data <= "0000000000";
                when x"1FC0" => data <= "0000000000";
                when x"1FC1" => data <= "0000000000";
                when x"1FC2" => data <= "0000000000";
                when x"1FC3" => data <= "0000000000";
                when x"1FC4" => data <= "0000000000";
                when x"1FC5" => data <= "0000000000";
                when x"1FC6" => data <= "0000000000";
                when x"1FC7" => data <= "0000000000";
                when x"1FC8" => data <= "0000000000";
                when x"1FC9" => data <= "0000000000";
                when x"1FCA" => data <= "0000000000";
                when x"1FCB" => data <= "0000000000";
                when x"1FCC" => data <= "0000000000";
                when x"1FCD" => data <= "0000000000";
                when x"1FCE" => data <= "0000000000";
                when x"1FCF" => data <= "0000000000";
                when x"1FD0" => data <= "0000000000";
                when x"1FD1" => data <= "0000000000";
                when x"1FD2" => data <= "0000000000";
                when x"1FD3" => data <= "0000000000";
                when x"1FD4" => data <= "0000000000";
                when x"1FD5" => data <= "0000000000";
                when x"1FD6" => data <= "0000000000";
                when x"1FD7" => data <= "0000000000";
                when x"1FD8" => data <= "0000000000";
                when x"1FD9" => data <= "0000000000";
                when x"1FDA" => data <= "0000000000";
                when x"1FDB" => data <= "0000000000";
                when x"1FDC" => data <= "0000000000";
                when x"1FDD" => data <= "0000000000";
                when x"1FDE" => data <= "0000000000";
                when x"1FDF" => data <= "0000000000";
                when x"1FE0" => data <= "0000000000";
                when x"1FE1" => data <= "0000000000";
                when x"1FE2" => data <= "0000000000";
                when x"1FE3" => data <= "0000000000";
                when x"1FE4" => data <= "0000000000";
                when x"1FE5" => data <= "0000000000";
                when x"1FE6" => data <= "0000000000";
                when x"1FE7" => data <= "0000000000";
                when x"1FE8" => data <= "0000000000";
                when x"1FE9" => data <= "0000000000";
                when x"1FEA" => data <= "0000000000";
                when x"1FEB" => data <= "0000000000";
                when x"1FEC" => data <= "0000000000";
                when x"1FED" => data <= "0000000000";
                when x"1FEE" => data <= "0000000000";
                when x"1FEF" => data <= "0000000000";
                when x"1FF0" => data <= "0000000000";
                when x"1FF1" => data <= "0000000000";
                when x"1FF2" => data <= "0000000000";
                when x"1FF3" => data <= "0000000000";
                when x"1FF4" => data <= "0000000000";
                when x"1FF5" => data <= "0000000000";
                when x"1FF6" => data <= "0000000000";
                when x"1FF7" => data <= "0000000000";
                when x"1FF8" => data <= "0000000000";
                when x"1FF9" => data <= "0000000000";
                when x"1FFA" => data <= "0000000000";
                when x"1FFB" => data <= "0000000000";
                when x"1FFC" => data <= "0000000000";
                when x"1FFD" => data <= "0000000000";
                when x"1FFE" => data <= "0000000000";
                when x"1FFF" => data <= "0000000000";
                when x"2000" => data <= "0000000000";
                when x"2001" => data <= "0000000000";
                when x"2002" => data <= "0000000000";
                when x"2003" => data <= "0000000000";
                when x"2004" => data <= "0000000000";
                when x"2005" => data <= "0000000000";
                when x"2006" => data <= "0000000000";
                when x"2007" => data <= "0000000000";
                when x"2008" => data <= "0000000000";
                when x"2009" => data <= "0000000000";
                when x"200A" => data <= "0000000000";
                when x"200B" => data <= "0000000000";
                when x"200C" => data <= "0000000000";
                when x"200D" => data <= "0000000000";
                when x"200E" => data <= "0000000000";
                when x"200F" => data <= "0000000000";
                when x"2010" => data <= "0000000000";
                when x"2011" => data <= "0000000000";
                when x"2012" => data <= "0000000000";
                when x"2013" => data <= "0000000000";
                when x"2014" => data <= "0000000000";
                when x"2015" => data <= "0000000000";
                when x"2016" => data <= "0000000000";
                when x"2017" => data <= "0000000000";
                when x"2018" => data <= "0000000000";
                when x"2019" => data <= "0000000000";
                when x"201A" => data <= "0000000000";
                when x"201B" => data <= "0000000000";
                when x"201C" => data <= "0000000000";
                when x"201D" => data <= "0000000000";
                when x"201E" => data <= "0000000000";
                when x"201F" => data <= "0000000000";
                when x"2020" => data <= "0000000000";
                when x"2021" => data <= "0000000000";
                when x"2022" => data <= "0000000000";
                when x"2023" => data <= "0000000000";
                when x"2024" => data <= "1111011011";
                when x"2025" => data <= "0000000000";
                when x"2026" => data <= "0000000000";
                when x"2027" => data <= "0000000000";
                when x"2028" => data <= "0000000000";
                when x"2029" => data <= "0000000000";
                when x"202A" => data <= "0000000000";
                when x"202B" => data <= "0000000000";
                when x"202C" => data <= "0000000000";
                when x"202D" => data <= "0000000000";
                when x"202E" => data <= "0000000000";
                when x"202F" => data <= "0000000000";
                when x"2030" => data <= "0000000000";
                when x"2031" => data <= "0000000000";
                when x"2032" => data <= "0000000000";
                when x"2033" => data <= "0000000000";
                when x"2034" => data <= "0000000000";
                when x"2035" => data <= "0000000000";
                when x"2036" => data <= "0000000000";
                when x"2037" => data <= "0000000000";
                when x"2038" => data <= "0000000000";
                when x"2039" => data <= "0000000000";
                when x"203A" => data <= "0000000000";
                when x"203B" => data <= "0000000000";
                when x"203C" => data <= "0000000000";
                when x"203D" => data <= "0000000000";
                when x"203E" => data <= "0000000000";
                when x"203F" => data <= "0000000000";
                when x"2040" => data <= "0000000000";
                when x"2041" => data <= "0000000000";
                when x"2042" => data <= "0000000000";
                when x"2043" => data <= "0000000000";
                when x"2044" => data <= "0000000000";
                when x"2045" => data <= "0000000000";
                when x"2046" => data <= "0000000000";
                when x"2047" => data <= "0000000000";
                when x"2048" => data <= "0000000000";
                when x"2049" => data <= "0000000000";
                when x"204A" => data <= "0000000000";
                when x"204B" => data <= "0000000000";
                when x"204C" => data <= "0000000000";
                when x"204D" => data <= "0000000000";
                when x"204E" => data <= "0000000000";
                when x"204F" => data <= "0000000000";
                when x"2050" => data <= "0000000000";
                when x"2051" => data <= "0111110111";
                when x"2052" => data <= "0000000000";
                when x"2053" => data <= "0000000000";
                when x"2054" => data <= "0000000000";
                when x"2055" => data <= "0000000000";
                when x"2056" => data <= "0000000000";
                when x"2057" => data <= "0000000000";
                when x"2058" => data <= "0000000000";
                when x"2059" => data <= "0000000000";
                when x"205A" => data <= "0000000000";
                when x"205B" => data <= "0000000000";
                when x"205C" => data <= "0000000000";
                when x"205D" => data <= "0000000000";
                when x"205E" => data <= "0000000000";
                when x"205F" => data <= "0000000000";
                when x"2060" => data <= "0000000000";
                when x"2061" => data <= "0000000000";
                when x"2062" => data <= "0000000000";
                when x"2063" => data <= "0000000000";
                when x"2064" => data <= "0000000000";
                when x"2065" => data <= "0000000000";
                when x"2066" => data <= "0000000000";
                when x"2067" => data <= "0000000000";
                when x"2068" => data <= "0000000000";
                when x"2069" => data <= "0000000000";
                when x"206A" => data <= "0000000000";
                when x"206B" => data <= "0000000000";
                when x"206C" => data <= "0000000000";
                when x"206D" => data <= "0000000000";
                when x"206E" => data <= "0000000000";
                when x"206F" => data <= "0000000000";
                when x"2070" => data <= "0000000000";
                when x"2071" => data <= "0000000000";
                when x"2072" => data <= "0000000000";
                when x"2073" => data <= "0000000000";
                when x"2074" => data <= "0000000000";
                when x"2075" => data <= "0000000000";
                when x"2076" => data <= "0000000000";
                when x"2077" => data <= "0000000000";
                when x"2078" => data <= "0000000000";
                when x"2079" => data <= "0000000000";
                when x"207A" => data <= "0000000000";
                when x"207B" => data <= "0000000000";
                when x"207C" => data <= "0000000000";
                when x"207D" => data <= "0000000000";
                when x"207E" => data <= "0000000000";
                when x"207F" => data <= "0000000000";
                when x"2080" => data <= "0000000000";
                when x"2081" => data <= "0000000000";
                when x"2082" => data <= "0000000000";
                when x"2083" => data <= "0000000000";
                when x"2084" => data <= "0000000000";
                when x"2085" => data <= "0000000000";
                when x"2086" => data <= "0000000000";
                when x"2087" => data <= "0000000000";
                when x"2088" => data <= "0000000000";
                when x"2089" => data <= "0000000000";
                when x"208A" => data <= "0000000000";
                when x"208B" => data <= "0000000000";
                when x"208C" => data <= "0000000000";
                when x"208D" => data <= "0000000000";
                when x"208E" => data <= "0000000000";
                when x"208F" => data <= "0000000000";
                when x"2090" => data <= "0000000000";
                when x"2091" => data <= "0000000000";
                when x"2092" => data <= "0000000000";
                when x"2093" => data <= "0000000000";
                when x"2094" => data <= "0000000000";
                when x"2095" => data <= "0000000000";
                when x"2096" => data <= "0000000000";
                when x"2097" => data <= "0000000000";
                when x"2098" => data <= "0000000000";
                when x"2099" => data <= "0000000000";
                when x"209A" => data <= "0000000000";
                when x"209B" => data <= "0000000000";
                when x"209C" => data <= "0000000000";
                when x"209D" => data <= "0000000000";
                when x"209E" => data <= "0000000000";
                when x"209F" => data <= "0000000000";
                when x"20A0" => data <= "0000000000";
                when x"20A1" => data <= "0000000000";
                when x"20A2" => data <= "0000000000";
                when x"20A3" => data <= "0000000000";
                when x"20A4" => data <= "0000000000";
                when x"20A5" => data <= "0000000000";
                when x"20A6" => data <= "0000000000";
                when x"20A7" => data <= "0000000000";
                when x"20A8" => data <= "0000000000";
                when x"20A9" => data <= "0000000000";
                when x"20AA" => data <= "0000000000";
                when x"20AB" => data <= "0000000000";
                when x"20AC" => data <= "0000000000";
                when x"20AD" => data <= "0000000000";
                when x"20AE" => data <= "0000000000";
                when x"20AF" => data <= "0000000000";
                when x"20B0" => data <= "0000000000";
                when x"20B1" => data <= "0000000000";
                when x"20B2" => data <= "0000000000";
                when x"20B3" => data <= "0000000000";
                when x"20B4" => data <= "0000000000";
                when x"20B5" => data <= "0000000000";
                when x"20B6" => data <= "0000000000";
                when x"20B7" => data <= "0000000000";
                when x"20B8" => data <= "0000000000";
                when x"20B9" => data <= "0000000000";
                when x"20BA" => data <= "0000000000";
                when x"20BB" => data <= "0000000000";
                when x"20BC" => data <= "0000000000";
                when x"20BD" => data <= "0000000000";
                when x"20BE" => data <= "0000000000";
                when x"20BF" => data <= "0000000000";
                when x"20C0" => data <= "0000000000";
                when x"20C1" => data <= "0000000000";
                when x"20C2" => data <= "0000000000";
                when x"20C3" => data <= "0000000000";
                when x"20C4" => data <= "0000000000";
                when x"20C5" => data <= "0000000000";
                when x"20C6" => data <= "0000000000";
                when x"20C7" => data <= "0000000000";
                when x"20C8" => data <= "0000000000";
                when x"20C9" => data <= "0000000000";
                when x"20CA" => data <= "0000000000";
                when x"20CB" => data <= "0000000000";
                when x"20CC" => data <= "0000000000";
                when x"20CD" => data <= "0000000000";
                when x"20CE" => data <= "0000000000";
                when x"20CF" => data <= "0000000000";
                when x"20D0" => data <= "0000000000";
                when x"20D1" => data <= "0000000000";
                when x"20D2" => data <= "0000000000";
                when x"20D3" => data <= "0000000000";
                when x"20D4" => data <= "0000000000";
                when x"20D5" => data <= "0000000000";
                when x"20D6" => data <= "0000000000";
                when x"20D7" => data <= "0000000000";
                when x"20D8" => data <= "0000000000";
                when x"20D9" => data <= "0000000000";
                when x"20DA" => data <= "0000000000";
                when x"20DB" => data <= "0000000000";
                when x"20DC" => data <= "0000000000";
                when x"20DD" => data <= "0000000000";
                when x"20DE" => data <= "0000000000";
                when x"20DF" => data <= "0000000000";
                when x"20E0" => data <= "0000000000";
                when x"20E1" => data <= "0000000000";
                when x"20E2" => data <= "0000000000";
                when x"20E3" => data <= "0000000000";
                when x"20E4" => data <= "0000000000";
                when x"20E5" => data <= "0000000000";
                when x"20E6" => data <= "0000000000";
                when x"20E7" => data <= "0000000000";
                when x"20E8" => data <= "0000000000";
                when x"20E9" => data <= "0000000000";
                when x"20EA" => data <= "0000000000";
                when x"20EB" => data <= "0000000000";
                when x"20EC" => data <= "0000000000";
                when x"20ED" => data <= "0000000000";
                when x"20EE" => data <= "0000000000";
                when x"20EF" => data <= "0000000000";
                when x"20F0" => data <= "0000000000";
                when x"20F1" => data <= "0000000000";
                when x"20F2" => data <= "0000000000";
                when x"20F3" => data <= "0000000000";
                when x"20F4" => data <= "0000000000";
                when x"20F5" => data <= "0000000000";
                when x"20F6" => data <= "0000000000";
                when x"20F7" => data <= "0000000000";
                when x"20F8" => data <= "0000000000";
                when x"20F9" => data <= "0000000000";
                when x"20FA" => data <= "0000000000";
                when x"20FB" => data <= "0000000000";
                when x"20FC" => data <= "0000000000";
                when x"20FD" => data <= "0000000000";
                when x"20FE" => data <= "0000000000";
                when x"20FF" => data <= "0000000000";
                when x"2100" => data <= "0000000000";
                when x"2101" => data <= "0000000000";
                when x"2102" => data <= "0000000000";
                when x"2103" => data <= "0000000000";
                when x"2104" => data <= "0000000000";
                when x"2105" => data <= "0000000000";
                when x"2106" => data <= "0000000000";
                when x"2107" => data <= "0000000000";
                when x"2108" => data <= "0000000000";
                when x"2109" => data <= "0000000000";
                when x"210A" => data <= "0000000000";
                when x"210B" => data <= "0000000000";
                when x"210C" => data <= "0000000000";
                when x"210D" => data <= "0000000000";
                when x"210E" => data <= "0000000000";
                when x"210F" => data <= "0000000000";
                when x"2110" => data <= "0000000000";
                when x"2111" => data <= "0000000000";
                when x"2112" => data <= "0000000000";
                when x"2113" => data <= "0000000000";
                when x"2114" => data <= "0000000000";
                when x"2115" => data <= "0000000000";
                when x"2116" => data <= "0000000000";
                when x"2117" => data <= "0000000000";
                when x"2118" => data <= "0000000000";
                when x"2119" => data <= "0000000000";
                when x"211A" => data <= "0000000000";
                when x"211B" => data <= "0000000000";
                when x"211C" => data <= "0000000000";
                when x"211D" => data <= "0000000000";
                when x"211E" => data <= "0000000000";
                when x"211F" => data <= "0000000000";
                when x"2120" => data <= "0000000000";
                when x"2121" => data <= "0000000000";
                when x"2122" => data <= "0000000000";
                when x"2123" => data <= "0000000000";
                when x"2124" => data <= "0000000000";
                when x"2125" => data <= "0000000000";
                when x"2126" => data <= "0000000000";
                when x"2127" => data <= "0000000000";
                when x"2128" => data <= "0000000000";
                when x"2129" => data <= "0000000000";
                when x"212A" => data <= "0000000000";
                when x"212B" => data <= "0000000000";
                when x"212C" => data <= "0000000000";
                when x"212D" => data <= "0000000000";
                when x"212E" => data <= "0000000000";
                when x"212F" => data <= "0000000000";
                when x"2130" => data <= "0000000000";
                when x"2131" => data <= "0000000000";
                when x"2132" => data <= "0000000000";
                when x"2133" => data <= "0000000000";
                when x"2134" => data <= "0000000000";
                when x"2135" => data <= "0000000000";
                when x"2136" => data <= "0000000000";
                when x"2137" => data <= "0000000000";
                when x"2138" => data <= "0000000000";
                when x"2139" => data <= "0000000000";
                when x"213A" => data <= "0000000000";
                when x"213B" => data <= "0000000000";
                when x"213C" => data <= "0000000000";
                when x"213D" => data <= "0000000000";
                when x"213E" => data <= "0000000000";
                when x"213F" => data <= "0000000000";
                when x"2140" => data <= "0000000000";
                when x"2141" => data <= "0000000000";
                when x"2142" => data <= "0000000000";
                when x"2143" => data <= "0000000000";
                when x"2144" => data <= "0000000000";
                when x"2145" => data <= "0000000000";
                when x"2146" => data <= "0000000000";
                when x"2147" => data <= "0000000000";
                when x"2148" => data <= "0000000000";
                when x"2149" => data <= "0000000000";
                when x"214A" => data <= "0000000000";
                when x"214B" => data <= "0000000000";
                when x"214C" => data <= "0000000000";
                when x"214D" => data <= "0000000000";
                when x"214E" => data <= "0000000000";
                when x"214F" => data <= "0000000000";
                when x"2150" => data <= "0000000000";
                when x"2151" => data <= "0000000000";
                when x"2152" => data <= "0000000000";
                when x"2153" => data <= "0000000000";
                when x"2154" => data <= "0000000000";
                when x"2155" => data <= "0000000000";
                when x"2156" => data <= "0000000000";
                when x"2157" => data <= "0000000000";
                when x"2158" => data <= "0000000000";
                when x"2159" => data <= "0000000000";
                when x"215A" => data <= "0000000000";
                when x"215B" => data <= "0000000000";
                when x"215C" => data <= "0000000000";
                when x"215D" => data <= "0000000000";
                when x"215E" => data <= "0000000000";
                when x"215F" => data <= "0000000000";
                when x"2160" => data <= "0000000000";
                when x"2161" => data <= "0000000000";
                when x"2162" => data <= "0000000000";
                when x"2163" => data <= "0000000000";
                when x"2164" => data <= "0000000000";
                when x"2165" => data <= "0000000000";
                when x"2166" => data <= "0000000000";
                when x"2167" => data <= "0000000000";
                when x"2168" => data <= "0000000000";
                when x"2169" => data <= "0000000000";
                when x"216A" => data <= "0000000000";
                when x"216B" => data <= "0000000000";
                when x"216C" => data <= "0000000000";
                when x"216D" => data <= "0000000000";
                when x"216E" => data <= "0000000000";
                when x"216F" => data <= "0000000000";
                when x"2170" => data <= "0000000000";
                when x"2171" => data <= "0000000000";
                when x"2172" => data <= "0000000000";
                when x"2173" => data <= "0000000000";
                when x"2174" => data <= "0000000000";
                when x"2175" => data <= "0000000000";
                when x"2176" => data <= "0000000000";
                when x"2177" => data <= "0000000000";
                when x"2178" => data <= "0000000000";
                when x"2179" => data <= "0000000000";
                when x"217A" => data <= "0000000000";
                when x"217B" => data <= "0000000000";
                when x"217C" => data <= "0000000000";
                when x"217D" => data <= "0000000000";
                when x"217E" => data <= "0000000000";
                when x"217F" => data <= "0000000000";
                when x"2180" => data <= "0000000000";
                when x"2181" => data <= "0000000000";
                when x"2182" => data <= "0000000000";
                when x"2183" => data <= "0000000000";
                when x"2184" => data <= "0000000000";
                when x"2185" => data <= "0000000000";
                when x"2186" => data <= "0111110111";
                when x"2187" => data <= "0000000000";
                when x"2188" => data <= "0000000000";
                when x"2189" => data <= "0000000000";
                when x"218A" => data <= "0000000000";
                when x"218B" => data <= "0000000000";
                when x"218C" => data <= "0000000000";
                when x"218D" => data <= "0000000000";
                when x"218E" => data <= "0000000000";
                when x"218F" => data <= "0000000000";
                when x"2190" => data <= "0000000000";
                when x"2191" => data <= "0000000000";
                when x"2192" => data <= "0000000000";
                when x"2193" => data <= "0000000000";
                when x"2194" => data <= "0000000000";
                when x"2195" => data <= "0000000000";
                when x"2196" => data <= "0000000000";
                when x"2197" => data <= "0000000000";
                when x"2198" => data <= "0000000000";
                when x"2199" => data <= "0000000000";
                when x"219A" => data <= "0000000000";
                when x"219B" => data <= "0000000000";
                when x"219C" => data <= "0000000000";
                when x"219D" => data <= "0000000000";
                when x"219E" => data <= "0000000000";
                when x"219F" => data <= "0000000000";
                when x"21A0" => data <= "0000000000";
                when x"21A1" => data <= "0000000000";
                when x"21A2" => data <= "0000000000";
                when x"21A3" => data <= "0000000000";
                when x"21A4" => data <= "0000000000";
                when x"21A5" => data <= "0000000000";
                when x"21A6" => data <= "0000000000";
                when x"21A7" => data <= "0000000000";
                when x"21A8" => data <= "0000000000";
                when x"21A9" => data <= "0000000000";
                when x"21AA" => data <= "0000000000";
                when x"21AB" => data <= "0000000000";
                when x"21AC" => data <= "0000000000";
                when x"21AD" => data <= "0000000000";
                when x"21AE" => data <= "0000000000";
                when x"21AF" => data <= "0000000000";
                when x"21B0" => data <= "0000000000";
                when x"21B1" => data <= "0000000000";
                when x"21B2" => data <= "0000000000";
                when x"21B3" => data <= "0000000000";
                when x"21B4" => data <= "0000000000";
                when x"21B5" => data <= "0000000000";
                when x"21B6" => data <= "0000000000";
                when x"21B7" => data <= "0000000000";
                when x"21B8" => data <= "0000000000";
                when x"21B9" => data <= "0000000000";
                when x"21BA" => data <= "0000000000";
                when x"21BB" => data <= "0000000000";
                when x"21BC" => data <= "0000000000";
                when x"21BD" => data <= "0000000000";
                when x"21BE" => data <= "0000000000";
                when x"21BF" => data <= "0000000000";
                when x"21C0" => data <= "0000000000";
                when x"21C1" => data <= "0000000000";
                when x"21C2" => data <= "0000000000";
                when x"21C3" => data <= "0000000000";
                when x"21C4" => data <= "0000000000";
                when x"21C5" => data <= "0000000000";
                when x"21C6" => data <= "0000000000";
                when x"21C7" => data <= "0000000000";
                when x"21C8" => data <= "0000000000";
                when x"21C9" => data <= "0000000000";
                when x"21CA" => data <= "0000000000";
                when x"21CB" => data <= "0000000000";
                when x"21CC" => data <= "0000000000";
                when x"21CD" => data <= "0000000000";
                when x"21CE" => data <= "0000000000";
                when x"21CF" => data <= "0000000000";
                when x"21D0" => data <= "0000000000";
                when x"21D1" => data <= "0000000000";
                when x"21D2" => data <= "0000000000";
                when x"21D3" => data <= "0000000000";
                when x"21D4" => data <= "0000000000";
                when x"21D5" => data <= "0000000000";
                when x"21D6" => data <= "0000000000";
                when x"21D7" => data <= "0000000000";
                when x"21D8" => data <= "0000000000";
                when x"21D9" => data <= "0000000000";
                when x"21DA" => data <= "0000000000";
                when x"21DB" => data <= "0000000000";
                when x"21DC" => data <= "0000000000";
                when x"21DD" => data <= "0000000000";
                when x"21DE" => data <= "0000000000";
                when x"21DF" => data <= "0000000000";
                when x"21E0" => data <= "0000000000";
                when x"21E1" => data <= "0000000000";
                when x"21E2" => data <= "0000000000";
                when x"21E3" => data <= "0000000000";
                when x"21E4" => data <= "0000000000";
                when x"21E5" => data <= "0000000000";
                when x"21E6" => data <= "1111011011";
                when x"21E7" => data <= "0000000000";
                when x"21E8" => data <= "0000000000";
                when x"21E9" => data <= "0000000000";
                when x"21EA" => data <= "0000000000";
                when x"21EB" => data <= "0000000000";
                when x"21EC" => data <= "0000000000";
                when x"21ED" => data <= "0000000000";
                when x"21EE" => data <= "0000000000";
                when x"21EF" => data <= "0000000000";
                when x"21F0" => data <= "0000000000";
                when x"21F1" => data <= "0000000000";
                when x"21F2" => data <= "0000000000";
                when x"21F3" => data <= "0000000000";
                when x"21F4" => data <= "0000000000";
                when x"21F5" => data <= "0000000000";
                when x"21F6" => data <= "0000000000";
                when x"21F7" => data <= "0000000000";
                when x"21F8" => data <= "0000000000";
                when x"21F9" => data <= "0000000000";
                when x"21FA" => data <= "0000000000";
                when x"21FB" => data <= "0000000000";
                when x"21FC" => data <= "0000000000";
                when x"21FD" => data <= "0000000000";
                when x"21FE" => data <= "0000000000";
                when x"21FF" => data <= "0000000000";
                when x"2200" => data <= "0000000000";
                when x"2201" => data <= "0000000000";
                when x"2202" => data <= "0000000000";
                when x"2203" => data <= "0000000000";
                when x"2204" => data <= "0000000000";
                when x"2205" => data <= "0000000000";
                when x"2206" => data <= "0000000000";
                when x"2207" => data <= "0000000000";
                when x"2208" => data <= "0000000000";
                when x"2209" => data <= "0000000000";
                when x"220A" => data <= "0000000000";
                when x"220B" => data <= "0000000000";
                when x"220C" => data <= "0000000000";
                when x"220D" => data <= "0000000000";
                when x"220E" => data <= "0000000000";
                when x"220F" => data <= "0000000000";
                when x"2210" => data <= "0000000000";
                when x"2211" => data <= "0000000000";
                when x"2212" => data <= "0000000000";
                when x"2213" => data <= "0000000000";
                when x"2214" => data <= "0000000000";
                when x"2215" => data <= "0000000000";
                when x"2216" => data <= "0000000000";
                when x"2217" => data <= "0000000000";
                when x"2218" => data <= "0000000000";
                when x"2219" => data <= "0000000000";
                when x"221A" => data <= "0000000000";
                when x"221B" => data <= "0000000000";
                when x"221C" => data <= "0000000000";
                when x"221D" => data <= "0000000000";
                when x"221E" => data <= "0000000000";
                when x"221F" => data <= "0000000000";
                when x"2220" => data <= "0111110111";
                when x"2221" => data <= "0000000000";
                when x"2222" => data <= "0000000000";
                when x"2223" => data <= "0111110111";
                when x"2224" => data <= "0000000000";
                when x"2225" => data <= "0000000000";
                when x"2226" => data <= "0000000000";
                when x"2227" => data <= "0000000000";
                when x"2228" => data <= "1101010000";
                when x"2229" => data <= "0000000000";
                when x"222A" => data <= "0000000000";
                when x"222B" => data <= "0000000000";
                when x"222C" => data <= "0000000000";
                when x"222D" => data <= "0000000000";
                when x"222E" => data <= "0000000000";
                when x"222F" => data <= "0000000000";
                when x"2230" => data <= "0000000000";
                when x"2231" => data <= "0000000000";
                when x"2232" => data <= "0000000000";
                when x"2233" => data <= "0000000000";
                when x"2234" => data <= "0000000000";
                when x"2235" => data <= "0000000000";
                when x"2236" => data <= "0000000000";
                when x"2237" => data <= "0000000000";
                when x"2238" => data <= "0000000000";
                when x"2239" => data <= "0000000000";
                when x"223A" => data <= "0000000000";
                when x"223B" => data <= "0000000000";
                when x"223C" => data <= "0000000000";
                when x"223D" => data <= "0000000000";
                when x"223E" => data <= "0000000000";
                when x"223F" => data <= "0000000000";
                when x"2240" => data <= "0000000000";
                when x"2241" => data <= "0000000000";
                when x"2242" => data <= "0000000000";
                when x"2243" => data <= "0000000000";
                when x"2244" => data <= "0000000000";
                when x"2245" => data <= "0000000000";
                when x"2246" => data <= "0000000000";
                when x"2247" => data <= "0000000000";
                when x"2248" => data <= "0000000000";
                when x"2249" => data <= "0000000000";
                when x"224A" => data <= "0000000000";
                when x"224B" => data <= "0000000000";
                when x"224C" => data <= "0000000000";
                when x"224D" => data <= "0000000000";
                when x"224E" => data <= "0000000000";
                when x"224F" => data <= "0000000000";
                when x"2250" => data <= "0000000000";
                when x"2251" => data <= "0000000000";
                when x"2252" => data <= "0000000000";
                when x"2253" => data <= "0000000000";
                when x"2254" => data <= "0000000000";
                when x"2255" => data <= "0000000000";
                when x"2256" => data <= "0000000000";
                when x"2257" => data <= "0000000000";
                when x"2258" => data <= "0000000000";
                when x"2259" => data <= "0000000000";
                when x"225A" => data <= "0000000000";
                when x"225B" => data <= "0000000000";
                when x"225C" => data <= "0000000000";
                when x"225D" => data <= "0000000000";
                when x"225E" => data <= "0000000000";
                when x"225F" => data <= "0000000000";
                when x"2260" => data <= "0000000000";
                when x"2261" => data <= "0000000000";
                when x"2262" => data <= "0000000000";
                when x"2263" => data <= "0000000000";
                when x"2264" => data <= "0000000000";
                when x"2265" => data <= "0000000000";
                when x"2266" => data <= "0000000000";
                when x"2267" => data <= "0000000000";
                when x"2268" => data <= "1101010000";
                when x"2269" => data <= "0000000000";
                when x"226A" => data <= "0000000000";
                when x"226B" => data <= "0000000000";
                when x"226C" => data <= "0000000000";
                when x"226D" => data <= "0000000000";
                when x"226E" => data <= "0000000000";
                when x"226F" => data <= "0000000000";
                when x"2270" => data <= "0000000000";
                when x"2271" => data <= "0000000000";
                when x"2272" => data <= "0000000000";
                when x"2273" => data <= "0000000000";
                when x"2274" => data <= "0000000000";
                when x"2275" => data <= "0000000000";
                when x"2276" => data <= "0000000000";
                when x"2277" => data <= "0000000000";
                when x"2278" => data <= "0000000000";
                when x"2279" => data <= "0000000000";
                when x"227A" => data <= "0000000000";
                when x"227B" => data <= "0000000000";
                when x"227C" => data <= "0000000000";
                when x"227D" => data <= "0000000000";
                when x"227E" => data <= "0000000000";
                when x"227F" => data <= "0000000000";
                when x"2280" => data <= "0000000000";
                when x"2281" => data <= "0000000000";
                when x"2282" => data <= "0000000000";
                when x"2283" => data <= "0000000000";
                when x"2284" => data <= "0000000000";
                when x"2285" => data <= "0000000000";
                when x"2286" => data <= "0000000000";
                when x"2287" => data <= "0000000000";
                when x"2288" => data <= "0000000000";
                when x"2289" => data <= "0000000000";
                when x"228A" => data <= "0000000000";
                when x"228B" => data <= "0000000000";
                when x"228C" => data <= "0000000000";
                when x"228D" => data <= "0000000000";
                when x"228E" => data <= "0000000000";
                when x"228F" => data <= "0000000000";
                when x"2290" => data <= "0000000000";
                when x"2291" => data <= "0000000000";
                when x"2292" => data <= "0000000000";
                when x"2293" => data <= "0000000000";
                when x"2294" => data <= "0000000000";
                when x"2295" => data <= "0000000000";
                when x"2296" => data <= "0000000000";
                when x"2297" => data <= "0000000000";
                when x"2298" => data <= "0000000000";
                when x"2299" => data <= "0000000000";
                when x"229A" => data <= "0000000000";
                when x"229B" => data <= "0000000000";
                when x"229C" => data <= "0000000000";
                when x"229D" => data <= "0000000000";
                when x"229E" => data <= "0000000000";
                when x"229F" => data <= "0000000000";
                when x"22A0" => data <= "0000000000";
                when x"22A1" => data <= "0000000000";
                when x"22A2" => data <= "0000000000";
                when x"22A3" => data <= "0000000000";
                when x"22A4" => data <= "0000000000";
                when x"22A5" => data <= "0000000000";
                when x"22A6" => data <= "0000000000";
                when x"22A7" => data <= "0000000000";
                when x"22A8" => data <= "0000000000";
                when x"22A9" => data <= "0000000000";
                when x"22AA" => data <= "0000000000";
                when x"22AB" => data <= "0000000000";
                when x"22AC" => data <= "0000000000";
                when x"22AD" => data <= "0000000000";
                when x"22AE" => data <= "0000000000";
                when x"22AF" => data <= "0000000000";
                when x"22B0" => data <= "0000000000";
                when x"22B1" => data <= "0000000000";
                when x"22B2" => data <= "0000000000";
                when x"22B3" => data <= "0000000000";
                when x"22B4" => data <= "0000000000";
                when x"22B5" => data <= "0000000000";
                when x"22B6" => data <= "0000000000";
                when x"22B7" => data <= "0000000000";
                when x"22B8" => data <= "0000000000";
                when x"22B9" => data <= "0000000000";
                when x"22BA" => data <= "0000000000";
                when x"22BB" => data <= "0000000000";
                when x"22BC" => data <= "0000000000";
                when x"22BD" => data <= "0000000000";
                when x"22BE" => data <= "0000000000";
                when x"22BF" => data <= "0000000000";
                when x"22C0" => data <= "0000000000";
                when x"22C1" => data <= "0000000000";
                when x"22C2" => data <= "0000000000";
                when x"22C3" => data <= "0000000000";
                when x"22C4" => data <= "0000000000";
                when x"22C5" => data <= "0000000000";
                when x"22C6" => data <= "0000000000";
                when x"22C7" => data <= "0000000000";
                when x"22C8" => data <= "0000000000";
                when x"22C9" => data <= "0000000000";
                when x"22CA" => data <= "0000000000";
                when x"22CB" => data <= "0000000000";
                when x"22CC" => data <= "0000000000";
                when x"22CD" => data <= "0000000000";
                when x"22CE" => data <= "0000000000";
                when x"22CF" => data <= "0000000000";
                when x"22D0" => data <= "0000000000";
                when x"22D1" => data <= "0000000000";
                when x"22D2" => data <= "0000000000";
                when x"22D3" => data <= "0000000000";
                when x"22D4" => data <= "0000000000";
                when x"22D5" => data <= "0000000000";
                when x"22D6" => data <= "0000000000";
                when x"22D7" => data <= "0000000000";
                when x"22D8" => data <= "0000000000";
                when x"22D9" => data <= "0000000000";
                when x"22DA" => data <= "0000000000";
                when x"22DB" => data <= "0000000000";
                when x"22DC" => data <= "0000000000";
                when x"22DD" => data <= "0000000000";
                when x"22DE" => data <= "0000000000";
                when x"22DF" => data <= "0000000000";
                when x"22E0" => data <= "0000000000";
                when x"22E1" => data <= "0000000000";
                when x"22E2" => data <= "0000000000";
                when x"22E3" => data <= "0000000000";
                when x"22E4" => data <= "0000000000";
                when x"22E5" => data <= "0000000000";
                when x"22E6" => data <= "0000000000";
                when x"22E7" => data <= "0000000000";
                when x"22E8" => data <= "0000000000";
                when x"22E9" => data <= "0000000000";
                when x"22EA" => data <= "0000000000";
                when x"22EB" => data <= "0000000000";
                when x"22EC" => data <= "0000000000";
                when x"22ED" => data <= "0000000000";
                when x"22EE" => data <= "0000000000";
                when x"22EF" => data <= "0000000000";
                when x"22F0" => data <= "0000000000";
                when x"22F1" => data <= "0000000000";
                when x"22F2" => data <= "0000000000";
                when x"22F3" => data <= "0000000000";
                when x"22F4" => data <= "0000000000";
                when x"22F5" => data <= "0000000000";
                when x"22F6" => data <= "0000000000";
                when x"22F7" => data <= "0000000000";
                when x"22F8" => data <= "0000000000";
                when x"22F9" => data <= "0000000000";
                when x"22FA" => data <= "0000000000";
                when x"22FB" => data <= "0000000000";
                when x"22FC" => data <= "0000000000";
                when x"22FD" => data <= "0000000000";
                when x"22FE" => data <= "0000000000";
                when x"22FF" => data <= "0000000000";
                when x"2300" => data <= "0000000000";
                when x"2301" => data <= "0000000000";
                when x"2302" => data <= "0000000000";
                when x"2303" => data <= "0000000000";
                when x"2304" => data <= "0000000000";
                when x"2305" => data <= "0000000000";
                when x"2306" => data <= "0000000000";
                when x"2307" => data <= "0000000000";
                when x"2308" => data <= "0000000000";
                when x"2309" => data <= "0000000000";
                when x"230A" => data <= "0000000000";
                when x"230B" => data <= "0000000000";
                when x"230C" => data <= "0000000000";
                when x"230D" => data <= "0000000000";
                when x"230E" => data <= "0000000000";
                when x"230F" => data <= "0000000000";
                when x"2310" => data <= "0000000000";
                when x"2311" => data <= "0000000000";
                when x"2312" => data <= "0000000000";
                when x"2313" => data <= "0000000000";
                when x"2314" => data <= "0000000000";
                when x"2315" => data <= "0000000000";
                when x"2316" => data <= "0000000000";
                when x"2317" => data <= "0000000000";
                when x"2318" => data <= "0000000000";
                when x"2319" => data <= "0000000000";
                when x"231A" => data <= "0000000000";
                when x"231B" => data <= "0000000000";
                when x"231C" => data <= "0000000000";
                when x"231D" => data <= "0000000000";
                when x"231E" => data <= "0000000000";
                when x"231F" => data <= "0000000000";
                when x"2320" => data <= "0000000000";
                when x"2321" => data <= "0000000000";
                when x"2322" => data <= "0000000000";
                when x"2323" => data <= "0000000000";
                when x"2324" => data <= "0000000000";
                when x"2325" => data <= "0000000000";
                when x"2326" => data <= "0000000000";
                when x"2327" => data <= "0000000000";
                when x"2328" => data <= "0000000000";
                when x"2329" => data <= "0000000000";
                when x"232A" => data <= "0000000000";
                when x"232B" => data <= "0000000000";
                when x"232C" => data <= "0000000000";
                when x"232D" => data <= "0000000000";
                when x"232E" => data <= "0000000000";
                when x"232F" => data <= "0000000000";
                when x"2330" => data <= "0000000000";
                when x"2331" => data <= "0000000000";
                when x"2332" => data <= "0000000000";
                when x"2333" => data <= "0000000000";
                when x"2334" => data <= "0000000000";
                when x"2335" => data <= "0000000000";
                when x"2336" => data <= "0000000000";
                when x"2337" => data <= "0000000000";
                when x"2338" => data <= "0000000000";
                when x"2339" => data <= "0000000000";
                when x"233A" => data <= "0000000000";
                when x"233B" => data <= "0000000000";
                when x"233C" => data <= "0000000000";
                when x"233D" => data <= "0000000000";
                when x"233E" => data <= "0000000000";
                when x"233F" => data <= "0000000000";
                when x"2340" => data <= "0000000000";
                when x"2341" => data <= "0000000000";
                when x"2342" => data <= "0000000000";
                when x"2343" => data <= "0000000000";
                when x"2344" => data <= "0000000000";
                when x"2345" => data <= "0000000000";
                when x"2346" => data <= "0000000000";
                when x"2347" => data <= "0000000000";
                when x"2348" => data <= "0000000000";
                when x"2349" => data <= "0000000000";
                when x"234A" => data <= "0000000000";
                when x"234B" => data <= "0000000000";
                when x"234C" => data <= "0000000000";
                when x"234D" => data <= "0000000000";
                when x"234E" => data <= "0000000000";
                when x"234F" => data <= "0000000000";
                when x"2350" => data <= "0000000000";
                when x"2351" => data <= "0000000000";
                when x"2352" => data <= "0000000000";
                when x"2353" => data <= "0000000000";
                when x"2354" => data <= "0000000000";
                when x"2355" => data <= "0000000000";
                when x"2356" => data <= "0000000000";
                when x"2357" => data <= "0111110111";
                when x"2358" => data <= "0000000000";
                when x"2359" => data <= "0000000000";
                when x"235A" => data <= "0000000000";
                when x"235B" => data <= "0000000000";
                when x"235C" => data <= "0000000000";
                when x"235D" => data <= "0000000000";
                when x"235E" => data <= "0000000000";
                when x"235F" => data <= "0000000000";
                when x"2360" => data <= "0000000000";
                when x"2361" => data <= "0000000000";
                when x"2362" => data <= "0000000000";
                when x"2363" => data <= "0000000000";
                when x"2364" => data <= "0000000000";
                when x"2365" => data <= "0000000000";
                when x"2366" => data <= "0000000000";
                when x"2367" => data <= "0000000000";
                when x"2368" => data <= "0000000000";
                when x"2369" => data <= "0000000000";
                when x"236A" => data <= "0000000000";
                when x"236B" => data <= "0000000000";
                when x"236C" => data <= "0000000000";
                when x"236D" => data <= "0000000000";
                when x"236E" => data <= "0000000000";
                when x"236F" => data <= "0000000000";
                when x"2370" => data <= "0000000000";
                when x"2371" => data <= "0000000000";
                when x"2372" => data <= "0000000000";
                when x"2373" => data <= "0000000000";
                when x"2374" => data <= "0000000000";
                when x"2375" => data <= "0000000000";
                when x"2376" => data <= "0000000000";
                when x"2377" => data <= "0000000000";
                when x"2378" => data <= "0000000000";
                when x"2379" => data <= "0000000000";
                when x"237A" => data <= "0000000000";
                when x"237B" => data <= "0000000000";
                when x"237C" => data <= "0000000000";
                when x"237D" => data <= "0000000000";
                when x"237E" => data <= "0000000000";
                when x"237F" => data <= "0000000000";
                when x"2380" => data <= "0000000000";
                when x"2381" => data <= "0000000000";
                when x"2382" => data <= "0000000000";
                when x"2383" => data <= "0000000000";
                when x"2384" => data <= "0000000000";
                when x"2385" => data <= "1100111010";
                when x"2386" => data <= "0000000000";
                when x"2387" => data <= "0000000000";
                when x"2388" => data <= "0000000000";
                when x"2389" => data <= "0000000000";
                when x"238A" => data <= "0000000000";
                when x"238B" => data <= "0000000000";
                when x"238C" => data <= "0000000000";
                when x"238D" => data <= "0000000000";
                when x"238E" => data <= "0000000000";
                when x"238F" => data <= "0000000000";
                when x"2390" => data <= "0000000000";
                when x"2391" => data <= "0000000000";
                when x"2392" => data <= "0000000000";
                when x"2393" => data <= "0000000000";
                when x"2394" => data <= "0000000000";
                when x"2395" => data <= "0000000000";
                when x"2396" => data <= "0000000000";
                when x"2397" => data <= "0000000000";
                when x"2398" => data <= "0000000000";
                when x"2399" => data <= "0000000000";
                when x"239A" => data <= "0000000000";
                when x"239B" => data <= "0000000000";
                when x"239C" => data <= "0000000000";
                when x"239D" => data <= "0000000000";
                when x"239E" => data <= "0000000000";
                when x"239F" => data <= "0000000000";
                when x"23A0" => data <= "0000000000";
                when x"23A1" => data <= "0000000000";
                when x"23A2" => data <= "0000000000";
                when x"23A3" => data <= "0000000000";
                when x"23A4" => data <= "0000000000";
                when x"23A5" => data <= "0000000000";
                when x"23A6" => data <= "0000000000";
                when x"23A7" => data <= "0000000000";
                when x"23A8" => data <= "0000000000";
                when x"23A9" => data <= "0000000000";
                when x"23AA" => data <= "0000000000";
                when x"23AB" => data <= "0000000000";
                when x"23AC" => data <= "0000000000";
                when x"23AD" => data <= "0000000000";
                when x"23AE" => data <= "0000000000";
                when x"23AF" => data <= "0000000000";
                when x"23B0" => data <= "0000000000";
                when x"23B1" => data <= "0000000000";
                when x"23B2" => data <= "0000000000";
                when x"23B3" => data <= "0000000000";
                when x"23B4" => data <= "0000000000";
                when x"23B5" => data <= "0000000000";
                when x"23B6" => data <= "0000000000";
                when x"23B7" => data <= "0000000000";
                when x"23B8" => data <= "0000000000";
                when x"23B9" => data <= "0000000000";
                when x"23BA" => data <= "0000000000";
                when x"23BB" => data <= "0000000000";
                when x"23BC" => data <= "0000000000";
                when x"23BD" => data <= "0000000000";
                when x"23BE" => data <= "0000000000";
                when x"23BF" => data <= "0000000000";
                when x"23C0" => data <= "0000000000";
                when x"23C1" => data <= "0000000000";
                when x"23C2" => data <= "0000000000";
                when x"23C3" => data <= "0000000000";
                when x"23C4" => data <= "0000000000";
                when x"23C5" => data <= "0000000000";
                when x"23C6" => data <= "0000000000";
                when x"23C7" => data <= "0000000000";
                when x"23C8" => data <= "0000000000";
                when x"23C9" => data <= "0000000000";
                when x"23CA" => data <= "0000000000";
                when x"23CB" => data <= "0000000000";
                when x"23CC" => data <= "0000000000";
                when x"23CD" => data <= "0000000000";
                when x"23CE" => data <= "0000000000";
                when x"23CF" => data <= "0000000000";
                when x"23D0" => data <= "0000000000";
                when x"23D1" => data <= "0000000000";
                when x"23D2" => data <= "0000000000";
                when x"23D3" => data <= "0000000000";
                when x"23D4" => data <= "0000000000";
                when x"23D5" => data <= "0000000000";
                when x"23D6" => data <= "0000000000";
                when x"23D7" => data <= "0000000000";
                when x"23D8" => data <= "0000000000";
                when x"23D9" => data <= "0000000000";
                when x"23DA" => data <= "0000000000";
                when x"23DB" => data <= "0000000000";
                when x"23DC" => data <= "0000000000";
                when x"23DD" => data <= "0000000000";
                when x"23DE" => data <= "0000000000";
                when x"23DF" => data <= "0000000000";
                when x"23E0" => data <= "0000000000";
                when x"23E1" => data <= "0000000000";
                when x"23E2" => data <= "0000000000";
                when x"23E3" => data <= "0000000000";
                when x"23E4" => data <= "0000000000";
                when x"23E5" => data <= "0000000000";
                when x"23E6" => data <= "0000000000";
                when x"23E7" => data <= "0000000000";
                when x"23E8" => data <= "0000000000";
                when x"23E9" => data <= "0000000000";
                when x"23EA" => data <= "0000000000";
                when x"23EB" => data <= "0000000000";
                when x"23EC" => data <= "0000000000";
                when x"23ED" => data <= "0000000000";
                when x"23EE" => data <= "0000000000";
                when x"23EF" => data <= "0000000000";
                when x"23F0" => data <= "0000000000";
                when x"23F1" => data <= "0000000000";
                when x"23F2" => data <= "0000000000";
                when x"23F3" => data <= "0000000000";
                when x"23F4" => data <= "0000000000";
                when x"23F5" => data <= "0000000000";
                when x"23F6" => data <= "0000000000";
                when x"23F7" => data <= "0000000000";
                when x"23F8" => data <= "0000000000";
                when x"23F9" => data <= "0000000000";
                when x"23FA" => data <= "0000000000";
                when x"23FB" => data <= "0000000000";
                when x"23FC" => data <= "0000000000";
                when x"23FD" => data <= "0000000000";
                when x"23FE" => data <= "0000000000";
                when x"23FF" => data <= "0000000000";
                when x"2400" => data <= "0000000000";
                when x"2401" => data <= "0000000000";
                when x"2402" => data <= "0000000000";
                when x"2403" => data <= "0000000000";
                when x"2404" => data <= "0000000000";
                when x"2405" => data <= "0000000000";
                when x"2406" => data <= "0000000000";
                when x"2407" => data <= "0000000000";
                when x"2408" => data <= "0000000000";
                when x"2409" => data <= "0000000000";
                when x"240A" => data <= "0000000000";
                when x"240B" => data <= "0000000000";
                when x"240C" => data <= "0000000000";
                when x"240D" => data <= "0000000000";
                when x"240E" => data <= "0000000000";
                when x"240F" => data <= "0000000000";
                when x"2410" => data <= "0000000000";
                when x"2411" => data <= "0000000000";
                when x"2412" => data <= "0000000000";
                when x"2413" => data <= "0000000000";
                when x"2414" => data <= "0000000000";
                when x"2415" => data <= "0000000000";
                when x"2416" => data <= "0000000000";
                when x"2417" => data <= "0000000000";
                when x"2418" => data <= "0000000000";
                when x"2419" => data <= "0000000000";
                when x"241A" => data <= "0000000000";
                when x"241B" => data <= "0000000000";
                when x"241C" => data <= "0000000000";
                when x"241D" => data <= "0000000000";
                when x"241E" => data <= "0000000000";
                when x"241F" => data <= "0000000000";
                when x"2420" => data <= "0000000000";
                when x"2421" => data <= "0000000000";
                when x"2422" => data <= "0000000000";
                when x"2423" => data <= "0000000000";
                when x"2424" => data <= "0000000000";
                when x"2425" => data <= "0000000000";
                when x"2426" => data <= "0000000000";
                when x"2427" => data <= "0000000000";
                when x"2428" => data <= "0000000000";
                when x"2429" => data <= "0000000000";
                when x"242A" => data <= "0000000000";
                when x"242B" => data <= "0000000000";
                when x"242C" => data <= "0000000000";
                when x"242D" => data <= "0000000000";
                when x"242E" => data <= "0000000000";
                when x"242F" => data <= "0000000000";
                when x"2430" => data <= "0000000000";
                when x"2431" => data <= "0000000000";
                when x"2432" => data <= "0000000000";
                when x"2433" => data <= "0000000000";
                when x"2434" => data <= "0000000000";
                when x"2435" => data <= "0000000000";
                when x"2436" => data <= "0000000000";
                when x"2437" => data <= "0000000000";
                when x"2438" => data <= "0000000000";
                when x"2439" => data <= "0000000000";
                when x"243A" => data <= "0000000000";
                when x"243B" => data <= "0000000000";
                when x"243C" => data <= "0000000000";
                when x"243D" => data <= "0000000000";
                when x"243E" => data <= "0000000000";
                when x"243F" => data <= "0000000000";
                when x"2440" => data <= "0000000000";
                when x"2441" => data <= "0000000000";
                when x"2442" => data <= "0000000000";
                when x"2443" => data <= "0000000000";
                when x"2444" => data <= "0000000000";
                when x"2445" => data <= "0000000000";
                when x"2446" => data <= "0000000000";
                when x"2447" => data <= "0000000000";
                when x"2448" => data <= "0000000000";
                when x"2449" => data <= "0000000000";
                when x"244A" => data <= "0000000000";
                when x"244B" => data <= "0000000000";
                when x"244C" => data <= "0000000000";
                when x"244D" => data <= "0000000000";
                when x"244E" => data <= "0000000000";
                when x"244F" => data <= "0000000000";
                when x"2450" => data <= "0000000000";
                when x"2451" => data <= "0000000000";
                when x"2452" => data <= "0000000000";
                when x"2453" => data <= "0000000000";
                when x"2454" => data <= "0000000000";
                when x"2455" => data <= "0000000000";
                when x"2456" => data <= "0000000000";
                when x"2457" => data <= "0000000000";
                when x"2458" => data <= "0000000000";
                when x"2459" => data <= "0000000000";
                when x"245A" => data <= "0000000000";
                when x"245B" => data <= "0000000000";
                when x"245C" => data <= "0000000000";
                when x"245D" => data <= "0000000000";
                when x"245E" => data <= "0000000000";
                when x"245F" => data <= "0000000000";
                when x"2460" => data <= "0000000000";
                when x"2461" => data <= "0000000000";
                when x"2462" => data <= "0000000000";
                when x"2463" => data <= "0000000000";
                when x"2464" => data <= "0000000000";
                when x"2465" => data <= "0000000000";
                when x"2466" => data <= "0000000000";
                when x"2467" => data <= "0000000000";
                when x"2468" => data <= "0000000000";
                when x"2469" => data <= "0000000000";
                when x"246A" => data <= "0000000000";
                when x"246B" => data <= "0000000000";
                when x"246C" => data <= "0000000000";
                when x"246D" => data <= "0000000000";
                when x"246E" => data <= "0000000000";
                when x"246F" => data <= "0000000000";
                when x"2470" => data <= "0000000000";
                when x"2471" => data <= "0000000000";
                when x"2472" => data <= "0000000000";
                when x"2473" => data <= "0000000000";
                when x"2474" => data <= "0000000000";
                when x"2475" => data <= "0000000000";
                when x"2476" => data <= "0110101000";
                when x"2477" => data <= "0000000000";
                when x"2478" => data <= "0000000000";
                when x"2479" => data <= "0000000000";
                when x"247A" => data <= "0000000000";
                when x"247B" => data <= "0000000000";
                when x"247C" => data <= "0000000000";
                when x"247D" => data <= "0000000000";
                when x"247E" => data <= "0000000000";
                when x"247F" => data <= "0000000000";
                when x"2480" => data <= "0000000000";
                when x"2481" => data <= "0000000000";
                when x"2482" => data <= "0000000000";
                when x"2483" => data <= "0000000000";
                when x"2484" => data <= "0000000000";
                when x"2485" => data <= "0000000000";
                when x"2486" => data <= "0000000000";
                when x"2487" => data <= "0000000000";
                when x"2488" => data <= "0000000000";
                when x"2489" => data <= "0000000000";
                when x"248A" => data <= "0000000000";
                when x"248B" => data <= "0000000000";
                when x"248C" => data <= "0000000000";
                when x"248D" => data <= "0000000000";
                when x"248E" => data <= "0000000000";
                when x"248F" => data <= "0000000000";
                when x"2490" => data <= "0000000000";
                when x"2491" => data <= "0000000000";
                when x"2492" => data <= "0000000000";
                when x"2493" => data <= "0000000000";
                when x"2494" => data <= "0000000000";
                when x"2495" => data <= "0000000000";
                when x"2496" => data <= "0000000000";
                when x"2497" => data <= "0000000000";
                when x"2498" => data <= "0000000000";
                when x"2499" => data <= "0000000000";
                when x"249A" => data <= "0000000000";
                when x"249B" => data <= "0000000000";
                when x"249C" => data <= "0000000000";
                when x"249D" => data <= "0000000000";
                when x"249E" => data <= "0000000000";
                when x"249F" => data <= "0000000000";
                when x"24A0" => data <= "0000000000";
                when x"24A1" => data <= "0000000000";
                when x"24A2" => data <= "0000000000";
                when x"24A3" => data <= "0000000000";
                when x"24A4" => data <= "0000000000";
                when x"24A5" => data <= "0000000000";
                when x"24A6" => data <= "0000000000";
                when x"24A7" => data <= "0000000000";
                when x"24A8" => data <= "0000000000";
                when x"24A9" => data <= "0000000000";
                when x"24AA" => data <= "0000000000";
                when x"24AB" => data <= "0000000000";
                when x"24AC" => data <= "0000000000";
                when x"24AD" => data <= "0000000000";
                when x"24AE" => data <= "0000000000";
                when x"24AF" => data <= "0000000000";
                when x"24B0" => data <= "0000000000";
                when x"24B1" => data <= "0000000000";
                when x"24B2" => data <= "0000000000";
                when x"24B3" => data <= "0000000000";
                when x"24B4" => data <= "0000000000";
                when x"24B5" => data <= "0000000000";
                when x"24B6" => data <= "0000000000";
                when x"24B7" => data <= "0000000000";
                when x"24B8" => data <= "0000000000";
                when x"24B9" => data <= "0000000000";
                when x"24BA" => data <= "0000000000";
                when x"24BB" => data <= "0000000000";
                when x"24BC" => data <= "0000000000";
                when x"24BD" => data <= "0000000000";
                when x"24BE" => data <= "0000000000";
                when x"24BF" => data <= "0000000000";
                when x"24C0" => data <= "0000000000";
                when x"24C1" => data <= "0000000000";
                when x"24C2" => data <= "0000000000";
                when x"24C3" => data <= "0000000000";
                when x"24C4" => data <= "0000000000";
                when x"24C5" => data <= "0000000000";
                when x"24C6" => data <= "0000000000";
                when x"24C7" => data <= "0000000000";
                when x"24C8" => data <= "0000000000";
                when x"24C9" => data <= "0000000000";
                when x"24CA" => data <= "0000000000";
                when x"24CB" => data <= "0000000000";
                when x"24CC" => data <= "0000000000";
                when x"24CD" => data <= "0000000000";
                when x"24CE" => data <= "0000000000";
                when x"24CF" => data <= "0000000000";
                when x"24D0" => data <= "0000000000";
                when x"24D1" => data <= "0000000000";
                when x"24D2" => data <= "0000000000";
                when x"24D3" => data <= "0000000000";
                when x"24D4" => data <= "0000000000";
                when x"24D5" => data <= "0000000000";
                when x"24D6" => data <= "0000000000";
                when x"24D7" => data <= "0000000000";
                when x"24D8" => data <= "0000000000";
                when x"24D9" => data <= "0000000000";
                when x"24DA" => data <= "0000000000";
                when x"24DB" => data <= "0000000000";
                when x"24DC" => data <= "0000000000";
                when x"24DD" => data <= "0000000000";
                when x"24DE" => data <= "0000000000";
                when x"24DF" => data <= "0000000000";
                when x"24E0" => data <= "0000000000";
                when x"24E1" => data <= "0000000000";
                when x"24E2" => data <= "0000000000";
                when x"24E3" => data <= "0000000000";
                when x"24E4" => data <= "0000000000";
                when x"24E5" => data <= "0000000000";
                when x"24E6" => data <= "0000000000";
                when x"24E7" => data <= "0000000000";
                when x"24E8" => data <= "0000000000";
                when x"24E9" => data <= "0000000000";
                when x"24EA" => data <= "0000000000";
                when x"24EB" => data <= "0000000000";
                when x"24EC" => data <= "0000000000";
                when x"24ED" => data <= "0000000000";
                when x"24EE" => data <= "0000000000";
                when x"24EF" => data <= "0000000000";
                when x"24F0" => data <= "0000000000";
                when x"24F1" => data <= "0000000000";
                when x"24F2" => data <= "0000000000";
                when x"24F3" => data <= "0000000000";
                when x"24F4" => data <= "0000000000";
                when x"24F5" => data <= "0000000000";
                when x"24F6" => data <= "0000000000";
                when x"24F7" => data <= "0000000000";
                when x"24F8" => data <= "0000000000";
                when x"24F9" => data <= "0000000000";
                when x"24FA" => data <= "0000000000";
                when x"24FB" => data <= "0000000000";
                when x"24FC" => data <= "0000000000";
                when x"24FD" => data <= "0000000000";
                when x"24FE" => data <= "0000000000";
                when x"24FF" => data <= "0000000000";
                when x"2500" => data <= "0000000000";
                when x"2501" => data <= "0000000000";
                when x"2502" => data <= "0000000000";
                when x"2503" => data <= "0000000000";
                when x"2504" => data <= "0000000000";
                when x"2505" => data <= "0000000000";
                when x"2506" => data <= "0000000000";
                when x"2507" => data <= "0000000000";
                when x"2508" => data <= "0000000000";
                when x"2509" => data <= "0000000000";
                when x"250A" => data <= "0000000000";
                when x"250B" => data <= "0000000000";
                when x"250C" => data <= "0000000000";
                when x"250D" => data <= "0000000000";
                when x"250E" => data <= "0000000000";
                when x"250F" => data <= "0000000000";
                when x"2510" => data <= "0000000000";
                when x"2511" => data <= "0000000000";
                when x"2512" => data <= "0000000000";
                when x"2513" => data <= "0000000000";
                when x"2514" => data <= "0000000000";
                when x"2515" => data <= "0000000000";
                when x"2516" => data <= "0000000000";
                when x"2517" => data <= "0000000000";
                when x"2518" => data <= "0000000000";
                when x"2519" => data <= "0000000000";
                when x"251A" => data <= "0000000000";
                when x"251B" => data <= "0000000000";
                when x"251C" => data <= "0000000000";
                when x"251D" => data <= "0000000000";
                when x"251E" => data <= "1001110011";
                when x"251F" => data <= "0000000000";
                when x"2520" => data <= "0000000000";
                when x"2521" => data <= "0000000000";
                when x"2522" => data <= "0000000000";
                when x"2523" => data <= "0000000000";
                when x"2524" => data <= "0000000000";
                when x"2525" => data <= "0000000000";
                when x"2526" => data <= "0000000000";
                when x"2527" => data <= "0000000000";
                when x"2528" => data <= "0000000000";
                when x"2529" => data <= "0000000000";
                when x"252A" => data <= "0000000000";
                when x"252B" => data <= "0000000000";
                when x"252C" => data <= "0000000000";
                when x"252D" => data <= "0000000000";
                when x"252E" => data <= "0000000000";
                when x"252F" => data <= "0000000000";
                when x"2530" => data <= "0000000000";
                when x"2531" => data <= "0000000000";
                when x"2532" => data <= "0000000000";
                when x"2533" => data <= "0000000000";
                when x"2534" => data <= "0000000000";
                when x"2535" => data <= "0000000000";
                when x"2536" => data <= "0000000000";
                when x"2537" => data <= "0000000000";
                when x"2538" => data <= "0000000000";
                when x"2539" => data <= "0000000000";
                when x"253A" => data <= "0000000000";
                when x"253B" => data <= "0000000000";
                when x"253C" => data <= "0000000000";
                when x"253D" => data <= "0000000000";
                when x"253E" => data <= "0000000000";
                when x"253F" => data <= "0000000000";
                when x"2540" => data <= "0000000000";
                when x"2541" => data <= "0000000000";
                when x"2542" => data <= "0000000000";
                when x"2543" => data <= "0000000000";
                when x"2544" => data <= "0000000000";
                when x"2545" => data <= "0000000000";
                when x"2546" => data <= "0000000000";
                when x"2547" => data <= "0000000000";
                when x"2548" => data <= "0000000000";
                when x"2549" => data <= "0000000000";
                when x"254A" => data <= "0000000000";
                when x"254B" => data <= "0000000000";
                when x"254C" => data <= "0000000000";
                when x"254D" => data <= "0000000000";
                when x"254E" => data <= "0000000000";
                when x"254F" => data <= "0000000000";
                when x"2550" => data <= "0000000000";
                when x"2551" => data <= "0000000000";
                when x"2552" => data <= "0000000000";
                when x"2553" => data <= "0000000000";
                when x"2554" => data <= "0000000000";
                when x"2555" => data <= "0000000000";
                when x"2556" => data <= "0000000000";
                when x"2557" => data <= "0000000000";
                when x"2558" => data <= "0000000000";
                when x"2559" => data <= "0000000000";
                when x"255A" => data <= "0000000000";
                when x"255B" => data <= "0000000000";
                when x"255C" => data <= "0000000000";
                when x"255D" => data <= "0000000000";
                when x"255E" => data <= "0000000000";
                when x"255F" => data <= "0000000000";
                when x"2560" => data <= "0000000000";
                when x"2561" => data <= "0000000000";
                when x"2562" => data <= "0000000000";
                when x"2563" => data <= "0000000000";
                when x"2564" => data <= "0000000000";
                when x"2565" => data <= "0000000000";
                when x"2566" => data <= "0000000000";
                when x"2567" => data <= "0000000000";
                when x"2568" => data <= "0000000000";
                when x"2569" => data <= "0000000000";
                when x"256A" => data <= "0000000000";
                when x"256B" => data <= "0000000000";
                when x"256C" => data <= "0000000000";
                when x"256D" => data <= "0000000000";
                when x"256E" => data <= "0000000000";
                when x"256F" => data <= "0000000000";
                when x"2570" => data <= "0000000000";
                when x"2571" => data <= "0000000000";
                when x"2572" => data <= "0000000000";
                when x"2573" => data <= "0000000000";
                when x"2574" => data <= "0000000000";
                when x"2575" => data <= "0111110111";
                when x"2576" => data <= "0000000000";
                when x"2577" => data <= "0000000000";
                when x"2578" => data <= "0000000000";
                when x"2579" => data <= "0000000000";
                when x"257A" => data <= "0000000000";
                when x"257B" => data <= "0000000000";
                when x"257C" => data <= "0000000000";
                when x"257D" => data <= "0000000000";
                when x"257E" => data <= "0000000000";
                when x"257F" => data <= "0000000000";
                when x"2580" => data <= "0000000000";
                when x"2581" => data <= "0000000000";
                when x"2582" => data <= "0000000000";
                when x"2583" => data <= "0000000000";
                when x"2584" => data <= "0000000000";
                when x"2585" => data <= "0000000000";
                when x"2586" => data <= "0000000000";
                when x"2587" => data <= "0000000000";
                when x"2588" => data <= "0000000000";
                when x"2589" => data <= "0000000000";
                when x"258A" => data <= "0000000000";
                when x"258B" => data <= "0000000000";
                when x"258C" => data <= "0000000000";
                when x"258D" => data <= "0000000000";
                when x"258E" => data <= "0000000000";
                when x"258F" => data <= "0000000000";
                when x"2590" => data <= "0000000000";
                when x"2591" => data <= "0000000000";
                when x"2592" => data <= "0000000000";
                when x"2593" => data <= "0000000000";
                when x"2594" => data <= "0000000000";
                when x"2595" => data <= "0000000000";
                when x"2596" => data <= "0000000000";
                when x"2597" => data <= "0000000000";
                when x"2598" => data <= "0000000000";
                when x"2599" => data <= "0000000000";
                when x"259A" => data <= "0000000000";
                when x"259B" => data <= "0000000000";
                when x"259C" => data <= "0000000000";
                when x"259D" => data <= "0000000000";
                when x"259E" => data <= "0000000000";
                when x"259F" => data <= "0000000000";
                when x"25A0" => data <= "0000000000";
                when x"25A1" => data <= "0000000000";
                when x"25A2" => data <= "0000000000";
                when x"25A3" => data <= "0000000000";
                when x"25A4" => data <= "0000000000";
                when x"25A5" => data <= "0000000000";
                when x"25A6" => data <= "0000000000";
                when x"25A7" => data <= "0000000000";
                when x"25A8" => data <= "0000000000";
                when x"25A9" => data <= "0000000000";
                when x"25AA" => data <= "0000000000";
                when x"25AB" => data <= "0000000000";
                when x"25AC" => data <= "0000000000";
                when x"25AD" => data <= "0000000000";
                when x"25AE" => data <= "0000000000";
                when x"25AF" => data <= "0000000000";
                when x"25B0" => data <= "0000000000";
                when x"25B1" => data <= "0000000000";
                when x"25B2" => data <= "0000000000";
                when x"25B3" => data <= "0000000000";
                when x"25B4" => data <= "0000000000";
                when x"25B5" => data <= "0000000000";
                when x"25B6" => data <= "0000000000";
                when x"25B7" => data <= "0000000000";
                when x"25B8" => data <= "0000000000";
                when x"25B9" => data <= "0000000000";
                when x"25BA" => data <= "0000000000";
                when x"25BB" => data <= "0000000000";
                when x"25BC" => data <= "0000000000";
                when x"25BD" => data <= "0000000000";
                when x"25BE" => data <= "0000000000";
                when x"25BF" => data <= "0000000000";
                when x"25C0" => data <= "0000000000";
                when x"25C1" => data <= "0000000000";
                when x"25C2" => data <= "0000000000";
                when x"25C3" => data <= "0000000000";
                when x"25C4" => data <= "0000000000";
                when x"25C5" => data <= "0000000000";
                when x"25C6" => data <= "0000000000";
                when x"25C7" => data <= "0000000000";
                when x"25C8" => data <= "0000000000";
                when x"25C9" => data <= "0000000000";
                when x"25CA" => data <= "0000000000";
                when x"25CB" => data <= "0000000000";
                when x"25CC" => data <= "0000000000";
                when x"25CD" => data <= "0000000000";
                when x"25CE" => data <= "0000000000";
                when x"25CF" => data <= "0000000000";
                when x"25D0" => data <= "0000000000";
                when x"25D1" => data <= "0000000000";
                when x"25D2" => data <= "0000000000";
                when x"25D3" => data <= "0000000000";
                when x"25D4" => data <= "0000000000";
                when x"25D5" => data <= "0000000000";
                when x"25D6" => data <= "0000000000";
                when x"25D7" => data <= "0000000000";
                when x"25D8" => data <= "0000000000";
                when x"25D9" => data <= "0000000000";
                when x"25DA" => data <= "0000000000";
                when x"25DB" => data <= "0000000000";
                when x"25DC" => data <= "0000000000";
                when x"25DD" => data <= "0000000000";
                when x"25DE" => data <= "0000000000";
                when x"25DF" => data <= "0000000000";
                when x"25E0" => data <= "0000000000";
                when x"25E1" => data <= "0000000000";
                when x"25E2" => data <= "0000000000";
                when x"25E3" => data <= "0000000000";
                when x"25E4" => data <= "0000000000";
                when x"25E5" => data <= "0000000000";
                when x"25E6" => data <= "0000000000";
                when x"25E7" => data <= "0000000000";
                when x"25E8" => data <= "0000000000";
                when x"25E9" => data <= "0000000000";
                when x"25EA" => data <= "0000000000";
                when x"25EB" => data <= "0000000000";
                when x"25EC" => data <= "0000000000";
                when x"25ED" => data <= "0000000000";
                when x"25EE" => data <= "0000000000";
                when x"25EF" => data <= "0000000000";
                when x"25F0" => data <= "0000000000";
                when x"25F1" => data <= "0000000000";
                when x"25F2" => data <= "0000000000";
                when x"25F3" => data <= "0000000000";
                when x"25F4" => data <= "0000000000";
                when x"25F5" => data <= "0000000000";
                when x"25F6" => data <= "0000000000";
                when x"25F7" => data <= "0000000000";
                when x"25F8" => data <= "0000000000";
                when x"25F9" => data <= "0000000000";
                when x"25FA" => data <= "0000000000";
                when x"25FB" => data <= "0000000000";
                when x"25FC" => data <= "0000000000";
                when x"25FD" => data <= "0000000000";
                when x"25FE" => data <= "0000000000";
                when x"25FF" => data <= "0000000000";
                when x"2600" => data <= "0000000000";
                when x"2601" => data <= "0000000000";
                when x"2602" => data <= "0000000000";
                when x"2603" => data <= "0000000000";
                when x"2604" => data <= "0111110111";
                when x"2605" => data <= "0000000000";
                when x"2606" => data <= "0000000000";
                when x"2607" => data <= "0000000000";
                when x"2608" => data <= "0000000000";
                when x"2609" => data <= "0000000000";
                when x"260A" => data <= "0000000000";
                when x"260B" => data <= "0000000000";
                when x"260C" => data <= "0000000000";
                when x"260D" => data <= "0000000000";
                when x"260E" => data <= "0000000000";
                when x"260F" => data <= "0000000000";
                when x"2610" => data <= "0000000000";
                when x"2611" => data <= "0000000000";
                when x"2612" => data <= "0000000000";
                when x"2613" => data <= "0000000000";
                when x"2614" => data <= "0000000000";
                when x"2615" => data <= "0000000000";
                when x"2616" => data <= "0000000000";
                when x"2617" => data <= "0000000000";
                when x"2618" => data <= "0000000000";
                when x"2619" => data <= "0000000000";
                when x"261A" => data <= "0000000000";
                when x"261B" => data <= "0000000000";
                when x"261C" => data <= "0000000000";
                when x"261D" => data <= "0000000000";
                when x"261E" => data <= "0000000000";
                when x"261F" => data <= "0000000000";
                when x"2620" => data <= "0000000000";
                when x"2621" => data <= "0000000000";
                when x"2622" => data <= "0000000000";
                when x"2623" => data <= "0000000000";
                when x"2624" => data <= "0000000000";
                when x"2625" => data <= "0000000000";
                when x"2626" => data <= "0000000000";
                when x"2627" => data <= "0000000000";
                when x"2628" => data <= "0000000000";
                when x"2629" => data <= "0000000000";
                when x"262A" => data <= "0000000000";
                when x"262B" => data <= "0000000000";
                when x"262C" => data <= "0000000000";
                when x"262D" => data <= "0000000000";
                when x"262E" => data <= "0000000000";
                when x"262F" => data <= "0000000000";
                when x"2630" => data <= "0000000000";
                when x"2631" => data <= "0000000000";
                when x"2632" => data <= "0000000000";
                when x"2633" => data <= "0000000000";
                when x"2634" => data <= "0000000000";
                when x"2635" => data <= "0000000000";
                when x"2636" => data <= "0000000000";
                when x"2637" => data <= "0000000000";
                when x"2638" => data <= "0000000000";
                when x"2639" => data <= "0000000000";
                when x"263A" => data <= "0000000000";
                when x"263B" => data <= "0000000000";
                when x"263C" => data <= "0000000000";
                when x"263D" => data <= "0000000000";
                when x"263E" => data <= "0000000000";
                when x"263F" => data <= "0000000000";
                when x"2640" => data <= "0000000000";
                when x"2641" => data <= "0000000000";
                when x"2642" => data <= "0000000000";
                when x"2643" => data <= "0000000000";
                when x"2644" => data <= "0000000000";
                when x"2645" => data <= "0000000000";
                when x"2646" => data <= "0000000000";
                when x"2647" => data <= "0000000000";
                when x"2648" => data <= "0000000000";
                when x"2649" => data <= "0000000000";
                when x"264A" => data <= "0000000000";
                when x"264B" => data <= "0000000000";
                when x"264C" => data <= "0000000000";
                when x"264D" => data <= "0000000000";
                when x"264E" => data <= "0000000000";
                when x"264F" => data <= "0000000000";
                when x"2650" => data <= "0000000000";
                when x"2651" => data <= "0000000000";
                when x"2652" => data <= "0000000000";
                when x"2653" => data <= "0000000000";
                when x"2654" => data <= "0000000000";
                when x"2655" => data <= "0000000000";
                when x"2656" => data <= "0000000000";
                when x"2657" => data <= "0000000000";
                when x"2658" => data <= "0000000000";
                when x"2659" => data <= "0000000000";
                when x"265A" => data <= "0000000000";
                when x"265B" => data <= "0000000000";
                when x"265C" => data <= "0000000000";
                when x"265D" => data <= "0000000000";
                when x"265E" => data <= "0000000000";
                when x"265F" => data <= "0000000000";
                when x"2660" => data <= "0000000000";
                when x"2661" => data <= "0000000000";
                when x"2662" => data <= "0000000000";
                when x"2663" => data <= "0000000000";
                when x"2664" => data <= "0000000000";
                when x"2665" => data <= "0000000000";
                when x"2666" => data <= "0000000000";
                when x"2667" => data <= "0000000000";
                when x"2668" => data <= "0000000000";
                when x"2669" => data <= "0000000000";
                when x"266A" => data <= "0000000000";
                when x"266B" => data <= "0000000000";
                when x"266C" => data <= "0000000000";
                when x"266D" => data <= "0000000000";
                when x"266E" => data <= "0000000000";
                when x"266F" => data <= "0000000000";
                when x"2670" => data <= "0000000000";
                when x"2671" => data <= "0111110111";
                when x"2672" => data <= "0000000000";
                when x"2673" => data <= "0000000000";
                when x"2674" => data <= "0000000000";
                when x"2675" => data <= "0000000000";
                when x"2676" => data <= "0000000000";
                when x"2677" => data <= "0000000000";
                when x"2678" => data <= "0000000000";
                when x"2679" => data <= "0000000000";
                when x"267A" => data <= "0000000000";
                when x"267B" => data <= "0000000000";
                when x"267C" => data <= "0000000000";
                when x"267D" => data <= "0000000000";
                when x"267E" => data <= "0000000000";
                when x"267F" => data <= "0000000000";
                when x"2680" => data <= "0000000000";
                when x"2681" => data <= "0000000000";
                when x"2682" => data <= "0000000000";
                when x"2683" => data <= "0000000000";
                when x"2684" => data <= "0000000000";
                when x"2685" => data <= "0000000000";
                when x"2686" => data <= "0000000000";
                when x"2687" => data <= "0000000000";
                when x"2688" => data <= "0000000000";
                when x"2689" => data <= "0000000000";
                when x"268A" => data <= "0000000000";
                when x"268B" => data <= "0000000000";
                when x"268C" => data <= "0000000000";
                when x"268D" => data <= "0000000000";
                when x"268E" => data <= "0000000000";
                when x"268F" => data <= "0000000000";
                when x"2690" => data <= "0000000000";
                when x"2691" => data <= "0000000000";
                when x"2692" => data <= "0000000000";
                when x"2693" => data <= "0000000000";
                when x"2694" => data <= "0000000000";
                when x"2695" => data <= "0000000000";
                when x"2696" => data <= "0000000000";
                when x"2697" => data <= "0000000000";
                when x"2698" => data <= "0000000000";
                when x"2699" => data <= "0000000000";
                when x"269A" => data <= "0000000000";
                when x"269B" => data <= "0000000000";
                when x"269C" => data <= "0000000000";
                when x"269D" => data <= "0000000000";
                when x"269E" => data <= "0000000000";
                when x"269F" => data <= "0000000000";
                when x"26A0" => data <= "0000000000";
                when x"26A1" => data <= "0000000000";
                when x"26A2" => data <= "0000000000";
                when x"26A3" => data <= "0000000000";
                when x"26A4" => data <= "0000000000";
                when x"26A5" => data <= "0000000000";
                when x"26A6" => data <= "0000000000";
                when x"26A7" => data <= "0000000000";
                when x"26A8" => data <= "0000000000";
                when x"26A9" => data <= "0000000000";
                when x"26AA" => data <= "0000000000";
                when x"26AB" => data <= "0000000000";
                when x"26AC" => data <= "0000000000";
                when x"26AD" => data <= "0000000000";
                when x"26AE" => data <= "0000000000";
                when x"26AF" => data <= "0000000000";
                when x"26B0" => data <= "0000000000";
                when x"26B1" => data <= "0000000000";
                when x"26B2" => data <= "0000000000";
                when x"26B3" => data <= "0000000000";
                when x"26B4" => data <= "0000000000";
                when x"26B5" => data <= "0000000000";
                when x"26B6" => data <= "0000000000";
                when x"26B7" => data <= "0000000000";
                when x"26B8" => data <= "0000000000";
                when x"26B9" => data <= "0000000000";
                when x"26BA" => data <= "0000000000";
                when x"26BB" => data <= "0000000000";
                when x"26BC" => data <= "0000000000";
                when x"26BD" => data <= "0000000000";
                when x"26BE" => data <= "0000000000";
                when x"26BF" => data <= "0000000000";
                when x"26C0" => data <= "0000000000";
                when x"26C1" => data <= "0000000000";
                when x"26C2" => data <= "0000000000";
                when x"26C3" => data <= "0000000000";
                when x"26C4" => data <= "0000000000";
                when x"26C5" => data <= "0000000000";
                when x"26C6" => data <= "0000000000";
                when x"26C7" => data <= "0000000000";
                when x"26C8" => data <= "0000000000";
                when x"26C9" => data <= "0000000000";
                when x"26CA" => data <= "0000000000";
                when x"26CB" => data <= "0000000000";
                when x"26CC" => data <= "0000000000";
                when x"26CD" => data <= "0000000000";
                when x"26CE" => data <= "0000000000";
                when x"26CF" => data <= "0000000000";
                when x"26D0" => data <= "0000000000";
                when x"26D1" => data <= "0000000000";
                when x"26D2" => data <= "0000000000";
                when x"26D3" => data <= "0000000000";
                when x"26D4" => data <= "0000000000";
                when x"26D5" => data <= "0000000000";
                when x"26D6" => data <= "0000000000";
                when x"26D7" => data <= "0000000000";
                when x"26D8" => data <= "0000000000";
                when x"26D9" => data <= "0000000000";
                when x"26DA" => data <= "0000000000";
                when x"26DB" => data <= "0000000000";
                when x"26DC" => data <= "0000000000";
                when x"26DD" => data <= "0000000000";
                when x"26DE" => data <= "0000000000";
                when x"26DF" => data <= "0000000000";
                when x"26E0" => data <= "0000000000";
                when x"26E1" => data <= "0000000000";
                when x"26E2" => data <= "0000000000";
                when x"26E3" => data <= "0000000000";
                when x"26E4" => data <= "0000000000";
                when x"26E5" => data <= "0000000000";
                when x"26E6" => data <= "0000000000";
                when x"26E7" => data <= "0000000000";
                when x"26E8" => data <= "0000000000";
                when x"26E9" => data <= "0000000000";
                when x"26EA" => data <= "0000000000";
                when x"26EB" => data <= "0000000000";
                when x"26EC" => data <= "0000000000";
                when x"26ED" => data <= "0000000000";
                when x"26EE" => data <= "0000000000";
                when x"26EF" => data <= "0000000000";
                when x"26F0" => data <= "0000000000";
                when x"26F1" => data <= "0000000000";
                when x"26F2" => data <= "0000000000";
                when x"26F3" => data <= "0000000000";
                when x"26F4" => data <= "0000000000";
                when x"26F5" => data <= "0000000000";
                when x"26F6" => data <= "0000000000";
                when x"26F7" => data <= "0000000000";
                when x"26F8" => data <= "0000000000";
                when x"26F9" => data <= "0000000000";
                when x"26FA" => data <= "0000000000";
                when x"26FB" => data <= "0000000000";
                when x"26FC" => data <= "0000000000";
                when x"26FD" => data <= "0000000000";
                when x"26FE" => data <= "0000000000";
                when x"26FF" => data <= "0000000000";
                when x"2700" => data <= "0000000000";
                when x"2701" => data <= "0000000000";
                when x"2702" => data <= "0000000000";
                when x"2703" => data <= "0000000000";
                when x"2704" => data <= "0000000000";
                when x"2705" => data <= "0000000000";
                when x"2706" => data <= "0000000000";
                when x"2707" => data <= "0000000000";
                when x"2708" => data <= "0000000000";
                when x"2709" => data <= "0000000000";
                when x"270A" => data <= "0000000000";
                when x"270B" => data <= "0000000000";
                when x"270C" => data <= "0000000000";
                when x"270D" => data <= "0000000000";
                when x"270E" => data <= "0000000000";
                when x"270F" => data <= "0000000000";
                when x"2710" => data <= "0000000000";
                when x"2711" => data <= "0000000000";
                when x"2712" => data <= "0000000000";
                when x"2713" => data <= "0000000000";
                when x"2714" => data <= "0000000000";
                when x"2715" => data <= "0000000000";
                when x"2716" => data <= "0000000000";
                when x"2717" => data <= "0000000000";
                when x"2718" => data <= "0000000000";
                when x"2719" => data <= "0000000000";
                when x"271A" => data <= "0000000000";
                when x"271B" => data <= "0000000000";
                when x"271C" => data <= "0000000000";
                when x"271D" => data <= "0000000000";
                when x"271E" => data <= "0000000000";
                when x"271F" => data <= "0000000000";
                when x"2720" => data <= "0000000000";
                when x"2721" => data <= "0000000000";
                when x"2722" => data <= "0000000000";
                when x"2723" => data <= "0000000000";
                when x"2724" => data <= "0000000000";
                when x"2725" => data <= "0000000000";
                when x"2726" => data <= "0000000000";
                when x"2727" => data <= "0000000000";
                when x"2728" => data <= "0000000000";
                when x"2729" => data <= "0000000000";
                when x"272A" => data <= "0000000000";
                when x"272B" => data <= "0000000000";
                when x"272C" => data <= "0000000000";
                when x"272D" => data <= "0000000000";
                when x"272E" => data <= "0000000000";
                when x"272F" => data <= "0000000000";
                when x"2730" => data <= "0000000000";
                when x"2731" => data <= "0000000000";
                when x"2732" => data <= "0000000000";
                when x"2733" => data <= "0000000000";
                when x"2734" => data <= "0000000000";
                when x"2735" => data <= "0000000000";
                when x"2736" => data <= "0000000000";
                when x"2737" => data <= "0000000000";
                when x"2738" => data <= "0000000000";
                when x"2739" => data <= "0000000000";
                when x"273A" => data <= "0000000000";
                when x"273B" => data <= "0000000000";
                when x"273C" => data <= "0000000000";
                when x"273D" => data <= "0000000000";
                when x"273E" => data <= "0000000000";
                when x"273F" => data <= "0000000000";
                when x"2740" => data <= "0000000000";
                when x"2741" => data <= "0000000000";
                when x"2742" => data <= "0000000000";
                when x"2743" => data <= "0000000000";
                when x"2744" => data <= "0000000000";
                when x"2745" => data <= "0000000000";
                when x"2746" => data <= "0000000000";
                when x"2747" => data <= "0000000000";
                when x"2748" => data <= "0000000000";
                when x"2749" => data <= "0000000000";
                when x"274A" => data <= "0000000000";
                when x"274B" => data <= "0000000000";
                when x"274C" => data <= "0000000000";
                when x"274D" => data <= "0000000000";
                when x"274E" => data <= "0000000000";
                when x"274F" => data <= "0000000000";
                when x"2750" => data <= "0000000000";
                when x"2751" => data <= "0000000000";
                when x"2752" => data <= "0000000000";
                when x"2753" => data <= "0000000000";
                when x"2754" => data <= "0000000000";
                when x"2755" => data <= "0000000000";
                when x"2756" => data <= "0000000000";
                when x"2757" => data <= "0000000000";
                when x"2758" => data <= "0000000000";
                when x"2759" => data <= "0000000000";
                when x"275A" => data <= "0000000000";
                when x"275B" => data <= "0000000000";
                when x"275C" => data <= "0000000000";
                when x"275D" => data <= "0000000000";
                when x"275E" => data <= "0000000000";
                when x"275F" => data <= "0000000000";
                when x"2760" => data <= "0000000000";
                when x"2761" => data <= "0000000000";
                when x"2762" => data <= "0000000000";
                when x"2763" => data <= "0000000000";
                when x"2764" => data <= "0000000000";
                when x"2765" => data <= "0000000000";
                when x"2766" => data <= "0000000000";
                when x"2767" => data <= "0000000000";
                when x"2768" => data <= "0000000000";
                when x"2769" => data <= "0000000000";
                when x"276A" => data <= "0000000000";
                when x"276B" => data <= "0000000000";
                when x"276C" => data <= "0000000000";
                when x"276D" => data <= "0000000000";
                when x"276E" => data <= "0000000000";
                when x"276F" => data <= "0000000000";
                when x"2770" => data <= "0000000000";
                when x"2771" => data <= "0000000000";
                when x"2772" => data <= "0000000000";
                when x"2773" => data <= "0000000000";
                when x"2774" => data <= "0000000000";
                when x"2775" => data <= "0000000000";
                when x"2776" => data <= "0000000000";
                when x"2777" => data <= "0000000000";
                when x"2778" => data <= "0000000000";
                when x"2779" => data <= "0000000000";
                when x"277A" => data <= "0000000000";
                when x"277B" => data <= "0000000000";
                when x"277C" => data <= "0000000000";
                when x"277D" => data <= "0000000000";
                when x"277E" => data <= "0000000000";
                when x"277F" => data <= "0000000000";
                when x"2780" => data <= "0000000000";
                when x"2781" => data <= "0000000000";
                when x"2782" => data <= "0000000000";
                when x"2783" => data <= "0000000000";
                when x"2784" => data <= "0000000000";
                when x"2785" => data <= "0000000000";
                when x"2786" => data <= "0000000000";
                when x"2787" => data <= "0000000000";
                when x"2788" => data <= "0000000000";
                when x"2789" => data <= "0000000000";
                when x"278A" => data <= "0000000000";
                when x"278B" => data <= "0000000000";
                when x"278C" => data <= "0000000000";
                when x"278D" => data <= "0000000000";
                when x"278E" => data <= "0000000000";
                when x"278F" => data <= "0000000000";
                when x"2790" => data <= "0000000000";
                when x"2791" => data <= "0000000000";
                when x"2792" => data <= "0000000000";
                when x"2793" => data <= "0000000000";
                when x"2794" => data <= "0000000000";
                when x"2795" => data <= "0000000000";
                when x"2796" => data <= "0000000000";
                when x"2797" => data <= "0000000000";
                when x"2798" => data <= "0000000000";
                when x"2799" => data <= "0000000000";
                when x"279A" => data <= "0000000000";
                when x"279B" => data <= "0000000000";
                when x"279C" => data <= "0000000000";
                when x"279D" => data <= "0000000000";
                when x"279E" => data <= "0000000000";
                when x"279F" => data <= "0000000000";
                when x"27A0" => data <= "0000000000";
                when x"27A1" => data <= "0000000000";
                when x"27A2" => data <= "0000000000";
                when x"27A3" => data <= "0000000000";
                when x"27A4" => data <= "0000000000";
                when x"27A5" => data <= "0000000000";
                when x"27A6" => data <= "0000000000";
                when x"27A7" => data <= "0000000000";
                when x"27A8" => data <= "0000000000";
                when x"27A9" => data <= "0000000000";
                when x"27AA" => data <= "0000000000";
                when x"27AB" => data <= "0000000000";
                when x"27AC" => data <= "0000000000";
                when x"27AD" => data <= "0000000000";
                when x"27AE" => data <= "0000000000";
                when x"27AF" => data <= "0000000000";
                when x"27B0" => data <= "0000000000";
                when x"27B1" => data <= "0000000000";
                when x"27B2" => data <= "0000000000";
                when x"27B3" => data <= "0000000000";
                when x"27B4" => data <= "0000000000";
                when x"27B5" => data <= "0000000000";
                when x"27B6" => data <= "0000000000";
                when x"27B7" => data <= "0000000000";
                when x"27B8" => data <= "0000000000";
                when x"27B9" => data <= "0000000000";
                when x"27BA" => data <= "0000000000";
                when x"27BB" => data <= "0000000000";
                when x"27BC" => data <= "0000000000";
                when x"27BD" => data <= "0000000000";
                when x"27BE" => data <= "0000000000";
                when x"27BF" => data <= "0000000000";
                when x"27C0" => data <= "0000000000";
                when x"27C1" => data <= "0000000000";
                when x"27C2" => data <= "0000000000";
                when x"27C3" => data <= "0000000000";
                when x"27C4" => data <= "0000000000";
                when x"27C5" => data <= "0000000000";
                when x"27C6" => data <= "0000000000";
                when x"27C7" => data <= "0000000000";
                when x"27C8" => data <= "0000000000";
                when x"27C9" => data <= "0000000000";
                when x"27CA" => data <= "0000000000";
                when x"27CB" => data <= "0000000000";
                when x"27CC" => data <= "0000000000";
                when x"27CD" => data <= "0000000000";
                when x"27CE" => data <= "0000000000";
                when x"27CF" => data <= "0000000000";
                when x"27D0" => data <= "0000000000";
                when x"27D1" => data <= "0000000000";
                when x"27D2" => data <= "0000000000";
                when x"27D3" => data <= "0000000000";
                when x"27D4" => data <= "0000000000";
                when x"27D5" => data <= "0000000000";
                when x"27D6" => data <= "0000000000";
                when x"27D7" => data <= "0000000000";
                when x"27D8" => data <= "0000000000";
                when x"27D9" => data <= "0000000000";
                when x"27DA" => data <= "0000000000";
                when x"27DB" => data <= "0000000000";
                when x"27DC" => data <= "0000000000";
                when x"27DD" => data <= "0000000000";
                when x"27DE" => data <= "0000000000";
                when x"27DF" => data <= "0000000000";
                when x"27E0" => data <= "0000000000";
                when x"27E1" => data <= "0000000000";
                when x"27E2" => data <= "0000000000";
                when x"27E3" => data <= "0000000000";
                when x"27E4" => data <= "0000000000";
                when x"27E5" => data <= "0000000000";
                when x"27E6" => data <= "0000000000";
                when x"27E7" => data <= "0000000000";
                when x"27E8" => data <= "0000000000";
                when x"27E9" => data <= "0000000000";
                when x"27EA" => data <= "0000000000";
                when x"27EB" => data <= "0000000000";
                when x"27EC" => data <= "0000000000";
                when x"27ED" => data <= "0000000000";
                when x"27EE" => data <= "0000000000";
                when x"27EF" => data <= "0000000000";
                when x"27F0" => data <= "0000000000";
                when x"27F1" => data <= "0000000000";
                when x"27F2" => data <= "0000000000";
                when x"27F3" => data <= "0000000000";
                when x"27F4" => data <= "0000000000";
                when x"27F5" => data <= "0000000000";
                when x"27F6" => data <= "0000000000";
                when x"27F7" => data <= "0000000000";
                when x"27F8" => data <= "0000000000";
                when x"27F9" => data <= "0000000000";
                when x"27FA" => data <= "0000000000";
                when x"27FB" => data <= "0000000000";
                when x"27FC" => data <= "0000000000";
                when x"27FD" => data <= "0000000000";
                when x"27FE" => data <= "0000000000";
                when x"27FF" => data <= "0000000000";
                when others => data <= (others => '0');
            end case;
        end if;
    end process;
end Behavioral;

------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity dic_mapper is
  generic ( WIDTH : integer := 8168 );
  port(
    data_in  : in  std_logic_vector(WIDTH-1 downto 0);
    data_out : out std_logic_vector(WIDTH-1 downto 0)
  );
end entity;

architecture Behavioral of dic_mapper is
begin
     data_out(0) <= data_in(0);
     data_out(1) <= data_in(1);
     data_out(2) <= data_in(2);
     data_out(3) <= data_in(3);
     data_out(4) <= data_in(4);
     data_out(5) <= data_in(5);
     data_out(6) <= data_in(6);
     data_out(7) <= data_in(7);
     data_out(8) <= data_in(8);
     data_out(9) <= data_in(9);
     data_out(10) <= data_in(10);
     data_out(11) <= data_in(11);
     data_out(12) <= data_in(12);
     data_out(13) <= data_in(13);
     data_out(14) <= data_in(14);
     data_out(15) <= data_in(15);
     data_out(16) <= data_in(16);
     data_out(17) <= data_in(17);
     data_out(18) <= data_in(18);
     data_out(19) <= data_in(19);
     data_out(20) <= data_in(20);
     data_out(21) <= data_in(21);
     data_out(22) <= data_in(22);
     data_out(23) <= data_in(23);
     data_out(24) <= data_in(24);
     data_out(25) <= data_in(25);
     data_out(26) <= data_in(26);
     data_out(27) <= data_in(27);
     data_out(28) <= data_in(28);
     data_out(29) <= data_in(29);
     data_out(30) <= data_in(30);
     data_out(31) <= data_in(31);
     data_out(32) <= data_in(32);
     data_out(33) <= data_in(33);
     data_out(34) <= data_in(34);
     data_out(35) <= data_in(35);
     data_out(36) <= data_in(36);
     data_out(37) <= data_in(37);
     data_out(38) <= data_in(38);
     data_out(39) <= data_in(39);
     data_out(40) <= data_in(40);
     data_out(41) <= data_in(41);
     data_out(42) <= data_in(42);
     data_out(43) <= data_in(43);
     data_out(44) <= data_in(44);
     data_out(45) <= data_in(45);
     data_out(46) <= data_in(46);
     data_out(47) <= data_in(47);
     data_out(48) <= data_in(48);
     data_out(49) <= data_in(49);
     data_out(50) <= data_in(50);
     data_out(51) <= data_in(51);
     data_out(52) <= data_in(52);
     data_out(53) <= data_in(53);
     data_out(54) <= data_in(54);
     data_out(55) <= data_in(55);
     data_out(56) <= data_in(56);
     data_out(57) <= data_in(57);
     data_out(58) <= data_in(58);
     data_out(59) <= data_in(59);
     data_out(60) <= data_in(60);
     data_out(61) <= data_in(61);
     data_out(62) <= data_in(62);
     data_out(63) <= data_in(63);
     data_out(64) <= data_in(64);
     data_out(65) <= data_in(65);
     data_out(66) <= data_in(66);
     data_out(67) <= data_in(67);
     data_out(68) <= data_in(68);
     data_out(69) <= data_in(69);
     data_out(70) <= data_in(70);
     data_out(71) <= data_in(71);
     data_out(72) <= data_in(72);
     data_out(73) <= data_in(73);
     data_out(74) <= data_in(74);
     data_out(75) <= data_in(75);
     data_out(76) <= data_in(76);
     data_out(77) <= data_in(77);
     data_out(78) <= data_in(78);
     data_out(79) <= data_in(79);
     data_out(80) <= data_in(80);
     data_out(81) <= data_in(81);
     data_out(82) <= data_in(82);
     data_out(83) <= data_in(83);
     data_out(84) <= data_in(84);
     data_out(85) <= data_in(85);
     data_out(86) <= data_in(86);
     data_out(87) <= data_in(87);
     data_out(88) <= data_in(88);
     data_out(89) <= data_in(89);
     data_out(90) <= data_in(90);
     data_out(91) <= data_in(91);
     data_out(92) <= data_in(92);
     data_out(93) <= data_in(93);
     data_out(94) <= data_in(94);
     data_out(95) <= data_in(95);
     data_out(96) <= data_in(96);
     data_out(97) <= data_in(97);
     data_out(98) <= data_in(98);
     data_out(99) <= data_in(99);
     data_out(100) <= data_in(100);
     data_out(101) <= data_in(101);
     data_out(102) <= data_in(102);
     data_out(103) <= data_in(103);
     data_out(104) <= data_in(104);
     data_out(105) <= data_in(105);
     data_out(106) <= data_in(106);
     data_out(107) <= data_in(107);
     data_out(108) <= data_in(108);
     data_out(109) <= data_in(109);
     data_out(110) <= data_in(110);
     data_out(111) <= data_in(111);
     data_out(112) <= data_in(112);
     data_out(113) <= data_in(113);
     data_out(114) <= data_in(114);
     data_out(115) <= data_in(115);
     data_out(116) <= data_in(116);
     data_out(117) <= data_in(117);
     data_out(118) <= data_in(118);
     data_out(119) <= data_in(119);
     data_out(120) <= data_in(120);
     data_out(121) <= data_in(121);
     data_out(122) <= data_in(122);
     data_out(123) <= data_in(123);
     data_out(124) <= data_in(124);
     data_out(125) <= data_in(125);
     data_out(126) <= data_in(126);
     data_out(127) <= data_in(127);
     data_out(128) <= data_in(128);
     data_out(129) <= data_in(129);
     data_out(130) <= data_in(130);
     data_out(131) <= data_in(131);
     data_out(132) <= data_in(132);
     data_out(133) <= data_in(133);
     data_out(134) <= data_in(134);
     data_out(135) <= data_in(135);
     data_out(136) <= data_in(136);
     data_out(137) <= data_in(137);
     data_out(138) <= data_in(138);
     data_out(139) <= data_in(139);
     data_out(140) <= data_in(140);
     data_out(141) <= data_in(141);
     data_out(142) <= data_in(142);
     data_out(143) <= data_in(143);
     data_out(144) <= data_in(144);
     data_out(145) <= data_in(145);
     data_out(146) <= data_in(146);
     data_out(147) <= data_in(147);
     data_out(148) <= data_in(148);
     data_out(149) <= data_in(149);
     data_out(150) <= data_in(150);
     data_out(151) <= data_in(151);
     data_out(152) <= data_in(152);
     data_out(153) <= data_in(153);
     data_out(154) <= data_in(154);
     data_out(155) <= data_in(155);
     data_out(156) <= data_in(156);
     data_out(157) <= data_in(157);
     data_out(158) <= data_in(158);
     data_out(159) <= data_in(159);
     data_out(160) <= data_in(160);
     data_out(161) <= data_in(161);
     data_out(162) <= data_in(162);
     data_out(163) <= data_in(163);
     data_out(164) <= data_in(164);
     data_out(165) <= data_in(165);
     data_out(166) <= data_in(166);
     data_out(167) <= data_in(167);
     data_out(168) <= data_in(168);
     data_out(169) <= data_in(169);
     data_out(170) <= data_in(170);
     data_out(171) <= data_in(171);
     data_out(172) <= data_in(172);
     data_out(173) <= data_in(173);
     data_out(174) <= data_in(174);
     data_out(175) <= data_in(175);
     data_out(176) <= data_in(176);
     data_out(177) <= data_in(177);
     data_out(178) <= data_in(178);
     data_out(179) <= data_in(179);
     data_out(180) <= data_in(180);
     data_out(181) <= data_in(181);
     data_out(182) <= data_in(182);
     data_out(183) <= data_in(183);
     data_out(184) <= data_in(184);
     data_out(185) <= data_in(185);
     data_out(186) <= data_in(186);
     data_out(187) <= data_in(187);
     data_out(188) <= data_in(188);
     data_out(189) <= data_in(189);
     data_out(190) <= data_in(190);
     data_out(191) <= data_in(191);
     data_out(192) <= data_in(192);
     data_out(193) <= data_in(193);
     data_out(194) <= data_in(194);
     data_out(195) <= data_in(195);
     data_out(196) <= data_in(196);
     data_out(197) <= data_in(197);
     data_out(198) <= data_in(198);
     data_out(199) <= data_in(199);
     data_out(200) <= data_in(200);
     data_out(201) <= data_in(201);
     data_out(202) <= data_in(202);
     data_out(203) <= data_in(203);
     data_out(204) <= data_in(204);
     data_out(205) <= data_in(205);
     data_out(206) <= data_in(206);
     data_out(207) <= data_in(207);
     data_out(208) <= data_in(208);
     data_out(209) <= data_in(209);
     data_out(210) <= data_in(210);
     data_out(211) <= data_in(211);
     data_out(212) <= data_in(212);
     data_out(213) <= data_in(213);
     data_out(214) <= data_in(214);
     data_out(215) <= data_in(215);
     data_out(216) <= data_in(216);
     data_out(217) <= data_in(217);
     data_out(218) <= data_in(218);
     data_out(219) <= data_in(219);
     data_out(220) <= data_in(220);
     data_out(221) <= data_in(221);
     data_out(222) <= data_in(222);
     data_out(223) <= data_in(223);
     data_out(224) <= data_in(224);
     data_out(225) <= data_in(225);
     data_out(226) <= data_in(226);
     data_out(227) <= data_in(227);
     data_out(228) <= data_in(228);
     data_out(229) <= data_in(229);
     data_out(230) <= data_in(230);
     data_out(231) <= data_in(231);
     data_out(232) <= data_in(232);
     data_out(233) <= data_in(233);
     data_out(234) <= data_in(234);
     data_out(235) <= data_in(235);
     data_out(236) <= data_in(236);
     data_out(237) <= data_in(237);
     data_out(238) <= data_in(238);
     data_out(239) <= data_in(239);
     data_out(240) <= data_in(246);
     data_out(241) <= data_in(248);
     data_out(242) <= data_in(250);
     data_out(243) <= data_in(251);
     data_out(244) <= data_in(252);
     data_out(245) <= data_in(258);
     data_out(246) <= data_in(259);
     data_out(247) <= data_in(262);
     data_out(248) <= data_in(265);
     data_out(249) <= data_in(266);
     data_out(250) <= data_in(277);
     data_out(251) <= data_in(279);
     data_out(252) <= data_in(281);
     data_out(253) <= data_in(284);
     data_out(254) <= data_in(294);
     data_out(255) <= data_in(299);
     data_out(256) <= data_in(305);
     data_out(257) <= data_in(307);
     data_out(258) <= data_in(313);
     data_out(259) <= data_in(318);
     data_out(260) <= data_in(323);
     data_out(261) <= data_in(324);
     data_out(262) <= data_in(325);
     data_out(263) <= data_in(327);
     data_out(264) <= data_in(329);
     data_out(265) <= data_in(330);
     data_out(266) <= data_in(332);
     data_out(267) <= data_in(336);
     data_out(268) <= data_in(343);
     data_out(269) <= data_in(344);
     data_out(270) <= data_in(345);
     data_out(271) <= data_in(353);
     data_out(272) <= data_in(354);
     data_out(273) <= data_in(355);
     data_out(274) <= data_in(359);
     data_out(275) <= data_in(360);
     data_out(276) <= data_in(367);
     data_out(277) <= data_in(369);
     data_out(278) <= data_in(370);
     data_out(279) <= data_in(371);
     data_out(280) <= data_in(381);
     data_out(281) <= data_in(384);
     data_out(282) <= data_in(388);
     data_out(283) <= data_in(389);
     data_out(284) <= data_in(393);
     data_out(285) <= data_in(394);
     data_out(286) <= data_in(396);
     data_out(287) <= data_in(399);
     data_out(288) <= data_in(400);
     data_out(289) <= data_in(405);
     data_out(290) <= data_in(406);
     data_out(291) <= data_in(408);
     data_out(292) <= data_in(409);
     data_out(293) <= data_in(411);
     data_out(294) <= data_in(412);
     data_out(295) <= data_in(413);
     data_out(296) <= data_in(419);
     data_out(297) <= data_in(420);
     data_out(298) <= data_in(423);
     data_out(299) <= data_in(426);
     data_out(300) <= data_in(429);
     data_out(301) <= data_in(432);
     data_out(302) <= data_in(433);
     data_out(303) <= data_in(434);
     data_out(304) <= data_in(435);
     data_out(305) <= data_in(439);
     data_out(306) <= data_in(440);
     data_out(307) <= data_in(446);
     data_out(308) <= data_in(449);
     data_out(309) <= data_in(450);
     data_out(310) <= data_in(456);
     data_out(311) <= data_in(458);
     data_out(312) <= data_in(459);
     data_out(313) <= data_in(461);
     data_out(314) <= data_in(462);
     data_out(315) <= data_in(463);
     data_out(316) <= data_in(465);
     data_out(317) <= data_in(467);
     data_out(318) <= data_in(469);
     data_out(319) <= data_in(470);
     data_out(320) <= data_in(471);
     data_out(321) <= data_in(474);
     data_out(322) <= data_in(477);
     data_out(323) <= data_in(478);
     data_out(324) <= data_in(485);
     data_out(325) <= data_in(486);
     data_out(326) <= data_in(488);
     data_out(327) <= data_in(489);
     data_out(328) <= data_in(492);
     data_out(329) <= data_in(495);
     data_out(330) <= data_in(500);
     data_out(331) <= data_in(504);
     data_out(332) <= data_in(505);
     data_out(333) <= data_in(507);
     data_out(334) <= data_in(509);
     data_out(335) <= data_in(510);
     data_out(336) <= data_in(511);
     data_out(337) <= data_in(513);
     data_out(338) <= data_in(516);
     data_out(339) <= data_in(520);
     data_out(340) <= data_in(521);
     data_out(341) <= data_in(522);
     data_out(342) <= data_in(533);
     data_out(343) <= data_in(537);
     data_out(344) <= data_in(538);
     data_out(345) <= data_in(539);
     data_out(346) <= data_in(542);
     data_out(347) <= data_in(544);
     data_out(348) <= data_in(545);
     data_out(349) <= data_in(546);
     data_out(350) <= data_in(547);
     data_out(351) <= data_in(548);
     data_out(352) <= data_in(549);
     data_out(353) <= data_in(551);
     data_out(354) <= data_in(553);
     data_out(355) <= data_in(554);
     data_out(356) <= data_in(555);
     data_out(357) <= data_in(559);
     data_out(358) <= data_in(560);
     data_out(359) <= data_in(563);
     data_out(360) <= data_in(570);
     data_out(361) <= data_in(571);
     data_out(362) <= data_in(572);
     data_out(363) <= data_in(574);
     data_out(364) <= data_in(576);
     data_out(365) <= data_in(577);
     data_out(366) <= data_in(578);
     data_out(367) <= data_in(579);
     data_out(368) <= data_in(580);
     data_out(369) <= data_in(582);
     data_out(370) <= data_in(583);
     data_out(371) <= data_in(585);
     data_out(372) <= data_in(586);
     data_out(373) <= data_in(588);
     data_out(374) <= data_in(589);
     data_out(375) <= data_in(590);
     data_out(376) <= data_in(595);
     data_out(377) <= data_in(596);
     data_out(378) <= data_in(598);
     data_out(379) <= data_in(599);
     data_out(380) <= data_in(601);
     data_out(381) <= data_in(605);
     data_out(382) <= data_in(606);
     data_out(383) <= data_in(607);
     data_out(384) <= data_in(608);
     data_out(385) <= data_in(612);
     data_out(386) <= data_in(614);
     data_out(387) <= data_in(615);
     data_out(388) <= data_in(619);
     data_out(389) <= data_in(621);
     data_out(390) <= data_in(624);
     data_out(391) <= data_in(626);
     data_out(392) <= data_in(629);
     data_out(393) <= data_in(631);
     data_out(394) <= data_in(632);
     data_out(395) <= data_in(633);
     data_out(396) <= data_in(636);
     data_out(397) <= data_in(637);
     data_out(398) <= data_in(643);
     data_out(399) <= data_in(647);
     data_out(400) <= data_in(648);
     data_out(401) <= data_in(649);
     data_out(402) <= data_in(653);
     data_out(403) <= data_in(658);
     data_out(404) <= data_in(659);
     data_out(405) <= data_in(660);
     data_out(406) <= data_in(661);
     data_out(407) <= data_in(668);
     data_out(408) <= data_in(670);
     data_out(409) <= data_in(672);
     data_out(410) <= data_in(673);
     data_out(411) <= data_in(674);
     data_out(412) <= data_in(679);
     data_out(413) <= data_in(681);
     data_out(414) <= data_in(682);
     data_out(415) <= data_in(685);
     data_out(416) <= data_in(687);
     data_out(417) <= data_in(692);
     data_out(418) <= data_in(694);
     data_out(419) <= data_in(695);
     data_out(420) <= data_in(697);
     data_out(421) <= data_in(698);
     data_out(422) <= data_in(699);
     data_out(423) <= data_in(700);
     data_out(424) <= data_in(708);
     data_out(425) <= data_in(711);
     data_out(426) <= data_in(713);
     data_out(427) <= data_in(714);
     data_out(428) <= data_in(715);
     data_out(429) <= data_in(722);
     data_out(430) <= data_in(725);
     data_out(431) <= data_in(726);
     data_out(432) <= data_in(727);
     data_out(433) <= data_in(728);
     data_out(434) <= data_in(734);
     data_out(435) <= data_in(735);
     data_out(436) <= data_in(738);
     data_out(437) <= data_in(739);
     data_out(438) <= data_in(741);
     data_out(439) <= data_in(743);
     data_out(440) <= data_in(749);
     data_out(441) <= data_in(752);
     data_out(442) <= data_in(753);
     data_out(443) <= data_in(754);
     data_out(444) <= data_in(757);
     data_out(445) <= data_in(758);
     data_out(446) <= data_in(759);
     data_out(447) <= data_in(760);
     data_out(448) <= data_in(761);
     data_out(449) <= data_in(762);
     data_out(450) <= data_in(763);
     data_out(451) <= data_in(768);
     data_out(452) <= data_in(770);
     data_out(453) <= data_in(778);
     data_out(454) <= data_in(782);
     data_out(455) <= data_in(784);
     data_out(456) <= data_in(785);
     data_out(457) <= data_in(786);
     data_out(458) <= data_in(789);
     data_out(459) <= data_in(797);
     data_out(460) <= data_in(798);
     data_out(461) <= data_in(799);
     data_out(462) <= data_in(801);
     data_out(463) <= data_in(803);
     data_out(464) <= data_in(804);
     data_out(465) <= data_in(805);
     data_out(466) <= data_in(808);
     data_out(467) <= data_in(814);
     data_out(468) <= data_in(817);
     data_out(469) <= data_in(818);
     data_out(470) <= data_in(820);
     data_out(471) <= data_in(821);
     data_out(472) <= data_in(825);
     data_out(473) <= data_in(829);
     data_out(474) <= data_in(831);
     data_out(475) <= data_in(835);
     data_out(476) <= data_in(836);
     data_out(477) <= data_in(839);
     data_out(478) <= data_in(840);
     data_out(479) <= data_in(842);
     data_out(480) <= data_in(843);
     data_out(481) <= data_in(845);
     data_out(482) <= data_in(849);
     data_out(483) <= data_in(858);
     data_out(484) <= data_in(863);
     data_out(485) <= data_in(864);
     data_out(486) <= data_in(865);
     data_out(487) <= data_in(868);
     data_out(488) <= data_in(872);
     data_out(489) <= data_in(874);
     data_out(490) <= data_in(876);
     data_out(491) <= data_in(878);
     data_out(492) <= data_in(882);
     data_out(493) <= data_in(884);
     data_out(494) <= data_in(885);
     data_out(495) <= data_in(886);
     data_out(496) <= data_in(888);
     data_out(497) <= data_in(894);
     data_out(498) <= data_in(897);
     data_out(499) <= data_in(898);
     data_out(500) <= data_in(899);
     data_out(501) <= data_in(900);
     data_out(502) <= data_in(920);
     data_out(503) <= data_in(921);
     data_out(504) <= data_in(924);
     data_out(505) <= data_in(925);
     data_out(506) <= data_in(926);
     data_out(507) <= data_in(927);
     data_out(508) <= data_in(928);
     data_out(509) <= data_in(929);
     data_out(510) <= data_in(930);
     data_out(511) <= data_in(935);
     data_out(512) <= data_in(939);
     data_out(513) <= data_in(942);
     data_out(514) <= data_in(943);
     data_out(515) <= data_in(948);
     data_out(516) <= data_in(949);
     data_out(517) <= data_in(950);
     data_out(518) <= data_in(953);
     data_out(519) <= data_in(964);
     data_out(520) <= data_in(965);
     data_out(521) <= data_in(966);
     data_out(522) <= data_in(967);
     data_out(523) <= data_in(968);
     data_out(524) <= data_in(970);
     data_out(525) <= data_in(971);
     data_out(526) <= data_in(973);
     data_out(527) <= data_in(977);
     data_out(528) <= data_in(980);
     data_out(529) <= data_in(982);
     data_out(530) <= data_in(984);
     data_out(531) <= data_in(985);
     data_out(532) <= data_in(986);
     data_out(533) <= data_in(989);
     data_out(534) <= data_in(993);
     data_out(535) <= data_in(996);
     data_out(536) <= data_in(1001);
     data_out(537) <= data_in(1002);
     data_out(538) <= data_in(1004);
     data_out(539) <= data_in(1005);
     data_out(540) <= data_in(1008);
     data_out(541) <= data_in(1014);
     data_out(542) <= data_in(1015);
     data_out(543) <= data_in(1016);
     data_out(544) <= data_in(1017);
     data_out(545) <= data_in(1019);
     data_out(546) <= data_in(1024);
     data_out(547) <= data_in(1027);
     data_out(548) <= data_in(1029);
     data_out(549) <= data_in(1032);
     data_out(550) <= data_in(1033);
     data_out(551) <= data_in(1036);
     data_out(552) <= data_in(1037);
     data_out(553) <= data_in(1041);
     data_out(554) <= data_in(1043);
     data_out(555) <= data_in(1045);
     data_out(556) <= data_in(1051);
     data_out(557) <= data_in(1054);
     data_out(558) <= data_in(1055);
     data_out(559) <= data_in(1057);
     data_out(560) <= data_in(1059);
     data_out(561) <= data_in(1061);
     data_out(562) <= data_in(1063);
     data_out(563) <= data_in(1064);
     data_out(564) <= data_in(1065);
     data_out(565) <= data_in(1067);
     data_out(566) <= data_in(1070);
     data_out(567) <= data_in(1071);
     data_out(568) <= data_in(1074);
     data_out(569) <= data_in(1075);
     data_out(570) <= data_in(1079);
     data_out(571) <= data_in(1080);
     data_out(572) <= data_in(1081);
     data_out(573) <= data_in(1083);
     data_out(574) <= data_in(1084);
     data_out(575) <= data_in(1086);
     data_out(576) <= data_in(1088);
     data_out(577) <= data_in(1089);
     data_out(578) <= data_in(1095);
     data_out(579) <= data_in(1096);
     data_out(580) <= data_in(1099);
     data_out(581) <= data_in(1100);
     data_out(582) <= data_in(1102);
     data_out(583) <= data_in(1103);
     data_out(584) <= data_in(1108);
     data_out(585) <= data_in(1109);
     data_out(586) <= data_in(1111);
     data_out(587) <= data_in(1112);
     data_out(588) <= data_in(1116);
     data_out(589) <= data_in(1119);
     data_out(590) <= data_in(1120);
     data_out(591) <= data_in(1121);
     data_out(592) <= data_in(1122);
     data_out(593) <= data_in(1140);
     data_out(594) <= data_in(1141);
     data_out(595) <= data_in(1148);
     data_out(596) <= data_in(1149);
     data_out(597) <= data_in(1152);
     data_out(598) <= data_in(1161);
     data_out(599) <= data_in(1168);
     data_out(600) <= data_in(1171);
     data_out(601) <= data_in(1172);
     data_out(602) <= data_in(1173);
     data_out(603) <= data_in(1174);
     data_out(604) <= data_in(1176);
     data_out(605) <= data_in(1178);
     data_out(606) <= data_in(1180);
     data_out(607) <= data_in(1183);
     data_out(608) <= data_in(1185);
     data_out(609) <= data_in(1187);
     data_out(610) <= data_in(1190);
     data_out(611) <= data_in(1191);
     data_out(612) <= data_in(1192);
     data_out(613) <= data_in(1193);
     data_out(614) <= data_in(1195);
     data_out(615) <= data_in(1198);
     data_out(616) <= data_in(1199);
     data_out(617) <= data_in(1203);
     data_out(618) <= data_in(1207);
     data_out(619) <= data_in(1208);
     data_out(620) <= data_in(1210);
     data_out(621) <= data_in(1211);
     data_out(622) <= data_in(1212);
     data_out(623) <= data_in(1213);
     data_out(624) <= data_in(1215);
     data_out(625) <= data_in(1216);
     data_out(626) <= data_in(1217);
     data_out(627) <= data_in(1218);
     data_out(628) <= data_in(1219);
     data_out(629) <= data_in(1220);
     data_out(630) <= data_in(1223);
     data_out(631) <= data_in(1224);
     data_out(632) <= data_in(1225);
     data_out(633) <= data_in(1227);
     data_out(634) <= data_in(1228);
     data_out(635) <= data_in(1229);
     data_out(636) <= data_in(1230);
     data_out(637) <= data_in(1232);
     data_out(638) <= data_in(1233);
     data_out(639) <= data_in(1237);
     data_out(640) <= data_in(1239);
     data_out(641) <= data_in(1242);
     data_out(642) <= data_in(1247);
     data_out(643) <= data_in(1252);
     data_out(644) <= data_in(1254);
     data_out(645) <= data_in(1255);
     data_out(646) <= data_in(1257);
     data_out(647) <= data_in(1258);
     data_out(648) <= data_in(1260);
     data_out(649) <= data_in(1262);
     data_out(650) <= data_in(1263);
     data_out(651) <= data_in(1267);
     data_out(652) <= data_in(1271);
     data_out(653) <= data_in(1273);
     data_out(654) <= data_in(1277);
     data_out(655) <= data_in(1279);
     data_out(656) <= data_in(1280);
     data_out(657) <= data_in(1283);
     data_out(658) <= data_in(1285);
     data_out(659) <= data_in(1287);
     data_out(660) <= data_in(1298);
     data_out(661) <= data_in(1302);
     data_out(662) <= data_in(1304);
     data_out(663) <= data_in(1305);
     data_out(664) <= data_in(1308);
     data_out(665) <= data_in(1309);
     data_out(666) <= data_in(1310);
     data_out(667) <= data_in(1313);
     data_out(668) <= data_in(1323);
     data_out(669) <= data_in(1326);
     data_out(670) <= data_in(1327);
     data_out(671) <= data_in(1328);
     data_out(672) <= data_in(1332);
     data_out(673) <= data_in(1333);
     data_out(674) <= data_in(1338);
     data_out(675) <= data_in(1344);
     data_out(676) <= data_in(1345);
     data_out(677) <= data_in(1347);
     data_out(678) <= data_in(1349);
     data_out(679) <= data_in(1354);
     data_out(680) <= data_in(1358);
     data_out(681) <= data_in(1360);
     data_out(682) <= data_in(1362);
     data_out(683) <= data_in(1363);
     data_out(684) <= data_in(1364);
     data_out(685) <= data_in(1365);
     data_out(686) <= data_in(1366);
     data_out(687) <= data_in(1369);
     data_out(688) <= data_in(1372);
     data_out(689) <= data_in(1378);
     data_out(690) <= data_in(1381);
     data_out(691) <= data_in(1384);
     data_out(692) <= data_in(1385);
     data_out(693) <= data_in(1386);
     data_out(694) <= data_in(1389);
     data_out(695) <= data_in(1390);
     data_out(696) <= data_in(1399);
     data_out(697) <= data_in(1401);
     data_out(698) <= data_in(1406);
     data_out(699) <= data_in(1407);
     data_out(700) <= data_in(1412);
     data_out(701) <= data_in(1414);
     data_out(702) <= data_in(1415);
     data_out(703) <= data_in(1422);
     data_out(704) <= data_in(1424);
     data_out(705) <= data_in(1425);
     data_out(706) <= data_in(1426);
     data_out(707) <= data_in(1428);
     data_out(708) <= data_in(1431);
     data_out(709) <= data_in(1439);
     data_out(710) <= data_in(1440);
     data_out(711) <= data_in(1445);
     data_out(712) <= data_in(1447);
     data_out(713) <= data_in(1450);
     data_out(714) <= data_in(1453);
     data_out(715) <= data_in(1457);
     data_out(716) <= data_in(1459);
     data_out(717) <= data_in(1460);
     data_out(718) <= data_in(1466);
     data_out(719) <= data_in(1468);
     data_out(720) <= data_in(1469);
     data_out(721) <= data_in(1470);
     data_out(722) <= data_in(1476);
     data_out(723) <= data_in(1478);
     data_out(724) <= data_in(1480);
     data_out(725) <= data_in(1483);
     data_out(726) <= data_in(1485);
     data_out(727) <= data_in(1486);
     data_out(728) <= data_in(1487);
     data_out(729) <= data_in(1489);
     data_out(730) <= data_in(1491);
     data_out(731) <= data_in(1497);
     data_out(732) <= data_in(1499);
     data_out(733) <= data_in(1501);
     data_out(734) <= data_in(1504);
     data_out(735) <= data_in(1506);
     data_out(736) <= data_in(1507);
     data_out(737) <= data_in(1508);
     data_out(738) <= data_in(1509);
     data_out(739) <= data_in(1510);
     data_out(740) <= data_in(1511);
     data_out(741) <= data_in(1512);
     data_out(742) <= data_in(1513);
     data_out(743) <= data_in(1515);
     data_out(744) <= data_in(1517);
     data_out(745) <= data_in(1518);
     data_out(746) <= data_in(1521);
     data_out(747) <= data_in(1524);
     data_out(748) <= data_in(1532);
     data_out(749) <= data_in(1533);
     data_out(750) <= data_in(1536);
     data_out(751) <= data_in(1537);
     data_out(752) <= data_in(1538);
     data_out(753) <= data_in(1541);
     data_out(754) <= data_in(1545);
     data_out(755) <= data_in(1546);
     data_out(756) <= data_in(1548);
     data_out(757) <= data_in(1551);
     data_out(758) <= data_in(1553);
     data_out(759) <= data_in(1555);
     data_out(760) <= data_in(1557);
     data_out(761) <= data_in(1561);
     data_out(762) <= data_in(1567);
     data_out(763) <= data_in(1569);
     data_out(764) <= data_in(1571);
     data_out(765) <= data_in(1572);
     data_out(766) <= data_in(1575);
     data_out(767) <= data_in(1578);
     data_out(768) <= data_in(1584);
     data_out(769) <= data_in(1586);
     data_out(770) <= data_in(1587);
     data_out(771) <= data_in(1589);
     data_out(772) <= data_in(1590);
     data_out(773) <= data_in(1592);
     data_out(774) <= data_in(1593);
     data_out(775) <= data_in(1594);
     data_out(776) <= data_in(1596);
     data_out(777) <= data_in(1598);
     data_out(778) <= data_in(1600);
     data_out(779) <= data_in(1603);
     data_out(780) <= data_in(1604);
     data_out(781) <= data_in(1606);
     data_out(782) <= data_in(1608);
     data_out(783) <= data_in(1611);
     data_out(784) <= data_in(1613);
     data_out(785) <= data_in(1614);
     data_out(786) <= data_in(1620);
     data_out(787) <= data_in(1622);
     data_out(788) <= data_in(1624);
     data_out(789) <= data_in(1626);
     data_out(790) <= data_in(1628);
     data_out(791) <= data_in(1634);
     data_out(792) <= data_in(1637);
     data_out(793) <= data_in(1638);
     data_out(794) <= data_in(1640);
     data_out(795) <= data_in(1641);
     data_out(796) <= data_in(1643);
     data_out(797) <= data_in(1645);
     data_out(798) <= data_in(1646);
     data_out(799) <= data_in(1651);
     data_out(800) <= data_in(1659);
     data_out(801) <= data_in(1660);
     data_out(802) <= data_in(1664);
     data_out(803) <= data_in(1667);
     data_out(804) <= data_in(1668);
     data_out(805) <= data_in(1670);
     data_out(806) <= data_in(1671);
     data_out(807) <= data_in(1674);
     data_out(808) <= data_in(1675);
     data_out(809) <= data_in(1676);
     data_out(810) <= data_in(1678);
     data_out(811) <= data_in(1681);
     data_out(812) <= data_in(1682);
     data_out(813) <= data_in(1684);
     data_out(814) <= data_in(1685);
     data_out(815) <= data_in(1686);
     data_out(816) <= data_in(1687);
     data_out(817) <= data_in(1688);
     data_out(818) <= data_in(1689);
     data_out(819) <= data_in(1695);
     data_out(820) <= data_in(1699);
     data_out(821) <= data_in(1700);
     data_out(822) <= data_in(1701);
     data_out(823) <= data_in(1703);
     data_out(824) <= data_in(1705);
     data_out(825) <= data_in(1711);
     data_out(826) <= data_in(1712);
     data_out(827) <= data_in(1713);
     data_out(828) <= data_in(1717);
     data_out(829) <= data_in(1719);
     data_out(830) <= data_in(1720);
     data_out(831) <= data_in(1721);
     data_out(832) <= data_in(1723);
     data_out(833) <= data_in(1725);
     data_out(834) <= data_in(1726);
     data_out(835) <= data_in(1727);
     data_out(836) <= data_in(1728);
     data_out(837) <= data_in(1729);
     data_out(838) <= data_in(1730);
     data_out(839) <= data_in(1731);
     data_out(840) <= data_in(1737);
     data_out(841) <= data_in(1741);
     data_out(842) <= data_in(1742);
     data_out(843) <= data_in(1743);
     data_out(844) <= data_in(1744);
     data_out(845) <= data_in(1747);
     data_out(846) <= data_in(1748);
     data_out(847) <= data_in(1754);
     data_out(848) <= data_in(1762);
     data_out(849) <= data_in(1763);
     data_out(850) <= data_in(1764);
     data_out(851) <= data_in(1766);
     data_out(852) <= data_in(1767);
     data_out(853) <= data_in(1768);
     data_out(854) <= data_in(1770);
     data_out(855) <= data_in(1773);
     data_out(856) <= data_in(1777);
     data_out(857) <= data_in(1779);
     data_out(858) <= data_in(1780);
     data_out(859) <= data_in(1781);
     data_out(860) <= data_in(1782);
     data_out(861) <= data_in(1783);
     data_out(862) <= data_in(1786);
     data_out(863) <= data_in(1788);
     data_out(864) <= data_in(1789);
     data_out(865) <= data_in(1790);
     data_out(866) <= data_in(1793);
     data_out(867) <= data_in(1795);
     data_out(868) <= data_in(1800);
     data_out(869) <= data_in(1804);
     data_out(870) <= data_in(1809);
     data_out(871) <= data_in(1812);
     data_out(872) <= data_in(1818);
     data_out(873) <= data_in(1820);
     data_out(874) <= data_in(1821);
     data_out(875) <= data_in(1824);
     data_out(876) <= data_in(1827);
     data_out(877) <= data_in(1828);
     data_out(878) <= data_in(1833);
     data_out(879) <= data_in(1836);
     data_out(880) <= data_in(1839);
     data_out(881) <= data_in(1841);
     data_out(882) <= data_in(1842);
     data_out(883) <= data_in(1844);
     data_out(884) <= data_in(1847);
     data_out(885) <= data_in(1848);
     data_out(886) <= data_in(1850);
     data_out(887) <= data_in(1853);
     data_out(888) <= data_in(1854);
     data_out(889) <= data_in(1855);
     data_out(890) <= data_in(1858);
     data_out(891) <= data_in(1859);
     data_out(892) <= data_in(1869);
     data_out(893) <= data_in(1872);
     data_out(894) <= data_in(1875);
     data_out(895) <= data_in(1876);
     data_out(896) <= data_in(1878);
     data_out(897) <= data_in(1879);
     data_out(898) <= data_in(1883);
     data_out(899) <= data_in(1885);
     data_out(900) <= data_in(1886);
     data_out(901) <= data_in(1887);
     data_out(902) <= data_in(1890);
     data_out(903) <= data_in(1891);
     data_out(904) <= data_in(1892);
     data_out(905) <= data_in(1893);
     data_out(906) <= data_in(1895);
     data_out(907) <= data_in(1896);
     data_out(908) <= data_in(1897);
     data_out(909) <= data_in(1898);
     data_out(910) <= data_in(1899);
     data_out(911) <= data_in(1902);
     data_out(912) <= data_in(1904);
     data_out(913) <= data_in(1906);
     data_out(914) <= data_in(1908);
     data_out(915) <= data_in(1911);
     data_out(916) <= data_in(1912);
     data_out(917) <= data_in(1913);
     data_out(918) <= data_in(1914);
     data_out(919) <= data_in(1915);
     data_out(920) <= data_in(1916);
     data_out(921) <= data_in(1917);
     data_out(922) <= data_in(1919);
     data_out(923) <= data_in(1922);
     data_out(924) <= data_in(1924);
     data_out(925) <= data_in(1925);
     data_out(926) <= data_in(1926);
     data_out(927) <= data_in(1930);
     data_out(928) <= data_in(1933);
     data_out(929) <= data_in(1937);
     data_out(930) <= data_in(1938);
     data_out(931) <= data_in(1939);
     data_out(932) <= data_in(1945);
     data_out(933) <= data_in(1947);
     data_out(934) <= data_in(1948);
     data_out(935) <= data_in(1955);
     data_out(936) <= data_in(1957);
     data_out(937) <= data_in(1959);
     data_out(938) <= data_in(1960);
     data_out(939) <= data_in(1961);
     data_out(940) <= data_in(1964);
     data_out(941) <= data_in(1966);
     data_out(942) <= data_in(1971);
     data_out(943) <= data_in(1974);
     data_out(944) <= data_in(1979);
     data_out(945) <= data_in(1980);
     data_out(946) <= data_in(1982);
     data_out(947) <= data_in(1984);
     data_out(948) <= data_in(1986);
     data_out(949) <= data_in(1987);
     data_out(950) <= data_in(1990);
     data_out(951) <= data_in(1992);
     data_out(952) <= data_in(1996);
     data_out(953) <= data_in(2000);
     data_out(954) <= data_in(2001);
     data_out(955) <= data_in(2006);
     data_out(956) <= data_in(2007);
     data_out(957) <= data_in(2010);
     data_out(958) <= data_in(2012);
     data_out(959) <= data_in(2018);
     data_out(960) <= data_in(2020);
     data_out(961) <= data_in(2021);
     data_out(962) <= data_in(2022);
     data_out(963) <= data_in(2026);
     data_out(964) <= data_in(2028);
     data_out(965) <= data_in(2034);
     data_out(966) <= data_in(2035);
     data_out(967) <= data_in(2036);
     data_out(968) <= data_in(2037);
     data_out(969) <= data_in(2038);
     data_out(970) <= data_in(2039);
     data_out(971) <= data_in(2040);
     data_out(972) <= data_in(2041);
     data_out(973) <= data_in(2049);
     data_out(974) <= data_in(2051);
     data_out(975) <= data_in(2053);
     data_out(976) <= data_in(2060);
     data_out(977) <= data_in(2062);
     data_out(978) <= data_in(2064);
     data_out(979) <= data_in(2066);
     data_out(980) <= data_in(2071);
     data_out(981) <= data_in(2073);
     data_out(982) <= data_in(2075);
     data_out(983) <= data_in(2076);
     data_out(984) <= data_in(2077);
     data_out(985) <= data_in(2079);
     data_out(986) <= data_in(2080);
     data_out(987) <= data_in(2081);
     data_out(988) <= data_in(2082);
     data_out(989) <= data_in(2085);
     data_out(990) <= data_in(2086);
     data_out(991) <= data_in(2087);
     data_out(992) <= data_in(2088);
     data_out(993) <= data_in(2089);
     data_out(994) <= data_in(2091);
     data_out(995) <= data_in(2093);
     data_out(996) <= data_in(2098);
     data_out(997) <= data_in(2099);
     data_out(998) <= data_in(2100);
     data_out(999) <= data_in(2101);
     data_out(1000) <= data_in(2102);
     data_out(1001) <= data_in(2105);
     data_out(1002) <= data_in(2106);
     data_out(1003) <= data_in(2108);
     data_out(1004) <= data_in(2118);
     data_out(1005) <= data_in(2121);
     data_out(1006) <= data_in(2123);
     data_out(1007) <= data_in(2129);
     data_out(1008) <= data_in(2131);
     data_out(1009) <= data_in(2133);
     data_out(1010) <= data_in(2134);
     data_out(1011) <= data_in(2135);
     data_out(1012) <= data_in(2136);
     data_out(1013) <= data_in(2139);
     data_out(1014) <= data_in(2140);
     data_out(1015) <= data_in(2141);
     data_out(1016) <= data_in(2143);
     data_out(1017) <= data_in(2146);
     data_out(1018) <= data_in(2148);
     data_out(1019) <= data_in(2150);
     data_out(1020) <= data_in(2152);
     data_out(1021) <= data_in(2153);
     data_out(1022) <= data_in(2154);
     data_out(1023) <= data_in(2158);
     data_out(1024) <= data_in(2163);
     data_out(1025) <= data_in(2165);
     data_out(1026) <= data_in(2170);
     data_out(1027) <= data_in(2173);
     data_out(1028) <= data_in(2174);
     data_out(1029) <= data_in(2175);
     data_out(1030) <= data_in(2177);
     data_out(1031) <= data_in(2180);
     data_out(1032) <= data_in(2183);
     data_out(1033) <= data_in(2184);
     data_out(1034) <= data_in(2185);
     data_out(1035) <= data_in(2186);
     data_out(1036) <= data_in(2187);
     data_out(1037) <= data_in(2189);
     data_out(1038) <= data_in(2191);
     data_out(1039) <= data_in(2195);
     data_out(1040) <= data_in(2200);
     data_out(1041) <= data_in(2213);
     data_out(1042) <= data_in(2217);
     data_out(1043) <= data_in(2218);
     data_out(1044) <= data_in(2221);
     data_out(1045) <= data_in(2224);
     data_out(1046) <= data_in(2228);
     data_out(1047) <= data_in(2231);
     data_out(1048) <= data_in(2234);
     data_out(1049) <= data_in(2235);
     data_out(1050) <= data_in(2236);
     data_out(1051) <= data_in(2237);
     data_out(1052) <= data_in(2238);
     data_out(1053) <= data_in(2241);
     data_out(1054) <= data_in(2242);
     data_out(1055) <= data_in(2243);
     data_out(1056) <= data_in(2244);
     data_out(1057) <= data_in(2247);
     data_out(1058) <= data_in(2248);
     data_out(1059) <= data_in(2252);
     data_out(1060) <= data_in(2255);
     data_out(1061) <= data_in(2264);
     data_out(1062) <= data_in(2265);
     data_out(1063) <= data_in(2266);
     data_out(1064) <= data_in(2267);
     data_out(1065) <= data_in(2268);
     data_out(1066) <= data_in(2270);
     data_out(1067) <= data_in(2272);
     data_out(1068) <= data_in(2273);
     data_out(1069) <= data_in(2275);
     data_out(1070) <= data_in(2277);
     data_out(1071) <= data_in(2279);
     data_out(1072) <= data_in(2281);
     data_out(1073) <= data_in(2283);
     data_out(1074) <= data_in(2285);
     data_out(1075) <= data_in(2287);
     data_out(1076) <= data_in(2289);
     data_out(1077) <= data_in(2290);
     data_out(1078) <= data_in(2291);
     data_out(1079) <= data_in(2294);
     data_out(1080) <= data_in(2296);
     data_out(1081) <= data_in(2299);
     data_out(1082) <= data_in(2305);
     data_out(1083) <= data_in(2306);
     data_out(1084) <= data_in(2312);
     data_out(1085) <= data_in(2313);
     data_out(1086) <= data_in(2314);
     data_out(1087) <= data_in(2315);
     data_out(1088) <= data_in(2318);
     data_out(1089) <= data_in(2322);
     data_out(1090) <= data_in(2323);
     data_out(1091) <= data_in(2324);
     data_out(1092) <= data_in(2326);
     data_out(1093) <= data_in(2328);
     data_out(1094) <= data_in(2329);
     data_out(1095) <= data_in(2332);
     data_out(1096) <= data_in(2333);
     data_out(1097) <= data_in(2338);
     data_out(1098) <= data_in(2341);
     data_out(1099) <= data_in(2344);
     data_out(1100) <= data_in(2351);
     data_out(1101) <= data_in(2353);
     data_out(1102) <= data_in(2355);
     data_out(1103) <= data_in(2358);
     data_out(1104) <= data_in(2359);
     data_out(1105) <= data_in(2362);
     data_out(1106) <= data_in(2365);
     data_out(1107) <= data_in(2366);
     data_out(1108) <= data_in(2371);
     data_out(1109) <= data_in(2372);
     data_out(1110) <= data_in(2379);
     data_out(1111) <= data_in(2385);
     data_out(1112) <= data_in(2386);
     data_out(1113) <= data_in(2389);
     data_out(1114) <= data_in(2390);
     data_out(1115) <= data_in(2391);
     data_out(1116) <= data_in(2394);
     data_out(1117) <= data_in(2395);
     data_out(1118) <= data_in(2396);
     data_out(1119) <= data_in(2397);
     data_out(1120) <= data_in(2399);
     data_out(1121) <= data_in(2404);
     data_out(1122) <= data_in(2406);
     data_out(1123) <= data_in(2407);
     data_out(1124) <= data_in(2409);
     data_out(1125) <= data_in(2410);
     data_out(1126) <= data_in(2411);
     data_out(1127) <= data_in(2414);
     data_out(1128) <= data_in(2418);
     data_out(1129) <= data_in(2421);
     data_out(1130) <= data_in(2427);
     data_out(1131) <= data_in(2429);
     data_out(1132) <= data_in(2430);
     data_out(1133) <= data_in(2433);
     data_out(1134) <= data_in(2434);
     data_out(1135) <= data_in(2437);
     data_out(1136) <= data_in(2438);
     data_out(1137) <= data_in(2440);
     data_out(1138) <= data_in(2441);
     data_out(1139) <= data_in(2444);
     data_out(1140) <= data_in(2448);
     data_out(1141) <= data_in(2449);
     data_out(1142) <= data_in(2454);
     data_out(1143) <= data_in(2455);
     data_out(1144) <= data_in(2457);
     data_out(1145) <= data_in(2458);
     data_out(1146) <= data_in(2459);
     data_out(1147) <= data_in(2460);
     data_out(1148) <= data_in(2463);
     data_out(1149) <= data_in(2467);
     data_out(1150) <= data_in(2468);
     data_out(1151) <= data_in(2473);
     data_out(1152) <= data_in(2490);
     data_out(1153) <= data_in(2496);
     data_out(1154) <= data_in(2497);
     data_out(1155) <= data_in(2502);
     data_out(1156) <= data_in(2503);
     data_out(1157) <= data_in(2504);
     data_out(1158) <= data_in(2507);
     data_out(1159) <= data_in(2508);
     data_out(1160) <= data_in(2514);
     data_out(1161) <= data_in(2515);
     data_out(1162) <= data_in(2516);
     data_out(1163) <= data_in(2518);
     data_out(1164) <= data_in(2520);
     data_out(1165) <= data_in(2521);
     data_out(1166) <= data_in(2522);
     data_out(1167) <= data_in(2523);
     data_out(1168) <= data_in(2524);
     data_out(1169) <= data_in(2529);
     data_out(1170) <= data_in(2532);
     data_out(1171) <= data_in(2533);
     data_out(1172) <= data_in(2534);
     data_out(1173) <= data_in(2536);
     data_out(1174) <= data_in(2537);
     data_out(1175) <= data_in(2538);
     data_out(1176) <= data_in(2541);
     data_out(1177) <= data_in(2542);
     data_out(1178) <= data_in(2544);
     data_out(1179) <= data_in(2546);
     data_out(1180) <= data_in(2547);
     data_out(1181) <= data_in(2548);
     data_out(1182) <= data_in(2549);
     data_out(1183) <= data_in(2550);
     data_out(1184) <= data_in(2553);
     data_out(1185) <= data_in(2555);
     data_out(1186) <= data_in(2559);
     data_out(1187) <= data_in(2561);
     data_out(1188) <= data_in(2562);
     data_out(1189) <= data_in(2570);
     data_out(1190) <= data_in(2573);
     data_out(1191) <= data_in(2574);
     data_out(1192) <= data_in(2575);
     data_out(1193) <= data_in(2576);
     data_out(1194) <= data_in(2580);
     data_out(1195) <= data_in(2581);
     data_out(1196) <= data_in(2582);
     data_out(1197) <= data_in(2583);
     data_out(1198) <= data_in(2585);
     data_out(1199) <= data_in(2589);
     data_out(1200) <= data_in(2595);
     data_out(1201) <= data_in(2596);
     data_out(1202) <= data_in(2601);
     data_out(1203) <= data_in(2607);
     data_out(1204) <= data_in(2608);
     data_out(1205) <= data_in(2611);
     data_out(1206) <= data_in(2612);
     data_out(1207) <= data_in(2614);
     data_out(1208) <= data_in(2615);
     data_out(1209) <= data_in(2617);
     data_out(1210) <= data_in(2621);
     data_out(1211) <= data_in(2622);
     data_out(1212) <= data_in(2624);
     data_out(1213) <= data_in(2625);
     data_out(1214) <= data_in(2626);
     data_out(1215) <= data_in(2629);
     data_out(1216) <= data_in(2632);
     data_out(1217) <= data_in(2634);
     data_out(1218) <= data_in(2635);
     data_out(1219) <= data_in(2638);
     data_out(1220) <= data_in(2640);
     data_out(1221) <= data_in(2642);
     data_out(1222) <= data_in(2643);
     data_out(1223) <= data_in(2646);
     data_out(1224) <= data_in(2647);
     data_out(1225) <= data_in(2651);
     data_out(1226) <= data_in(2653);
     data_out(1227) <= data_in(2654);
     data_out(1228) <= data_in(2655);
     data_out(1229) <= data_in(2660);
     data_out(1230) <= data_in(2661);
     data_out(1231) <= data_in(2663);
     data_out(1232) <= data_in(2670);
     data_out(1233) <= data_in(2672);
     data_out(1234) <= data_in(2674);
     data_out(1235) <= data_in(2676);
     data_out(1236) <= data_in(2677);
     data_out(1237) <= data_in(2678);
     data_out(1238) <= data_in(2679);
     data_out(1239) <= data_in(2682);
     data_out(1240) <= data_in(2683);
     data_out(1241) <= data_in(2684);
     data_out(1242) <= data_in(2686);
     data_out(1243) <= data_in(2691);
     data_out(1244) <= data_in(2696);
     data_out(1245) <= data_in(2698);
     data_out(1246) <= data_in(2699);
     data_out(1247) <= data_in(2703);
     data_out(1248) <= data_in(2705);
     data_out(1249) <= data_in(2713);
     data_out(1250) <= data_in(2714);
     data_out(1251) <= data_in(2715);
     data_out(1252) <= data_in(2716);
     data_out(1253) <= data_in(2717);
     data_out(1254) <= data_in(2721);
     data_out(1255) <= data_in(2724);
     data_out(1256) <= data_in(2726);
     data_out(1257) <= data_in(2731);
     data_out(1258) <= data_in(2743);
     data_out(1259) <= data_in(2746);
     data_out(1260) <= data_in(2748);
     data_out(1261) <= data_in(2750);
     data_out(1262) <= data_in(2751);
     data_out(1263) <= data_in(2753);
     data_out(1264) <= data_in(2755);
     data_out(1265) <= data_in(2760);
     data_out(1266) <= data_in(2761);
     data_out(1267) <= data_in(2762);
     data_out(1268) <= data_in(2765);
     data_out(1269) <= data_in(2770);
     data_out(1270) <= data_in(2771);
     data_out(1271) <= data_in(2774);
     data_out(1272) <= data_in(2776);
     data_out(1273) <= data_in(2778);
     data_out(1274) <= data_in(2779);
     data_out(1275) <= data_in(2780);
     data_out(1276) <= data_in(2782);
     data_out(1277) <= data_in(2784);
     data_out(1278) <= data_in(2786);
     data_out(1279) <= data_in(2787);
     data_out(1280) <= data_in(2796);
     data_out(1281) <= data_in(2803);
     data_out(1282) <= data_in(2804);
     data_out(1283) <= data_in(2805);
     data_out(1284) <= data_in(2808);
     data_out(1285) <= data_in(2809);
     data_out(1286) <= data_in(2811);
     data_out(1287) <= data_in(2812);
     data_out(1288) <= data_in(2814);
     data_out(1289) <= data_in(2816);
     data_out(1290) <= data_in(2822);
     data_out(1291) <= data_in(2824);
     data_out(1292) <= data_in(2829);
     data_out(1293) <= data_in(2831);
     data_out(1294) <= data_in(2832);
     data_out(1295) <= data_in(2837);
     data_out(1296) <= data_in(2841);
     data_out(1297) <= data_in(2843);
     data_out(1298) <= data_in(2844);
     data_out(1299) <= data_in(2848);
     data_out(1300) <= data_in(2850);
     data_out(1301) <= data_in(2852);
     data_out(1302) <= data_in(2853);
     data_out(1303) <= data_in(2855);
     data_out(1304) <= data_in(2856);
     data_out(1305) <= data_in(2860);
     data_out(1306) <= data_in(2862);
     data_out(1307) <= data_in(2863);
     data_out(1308) <= data_in(2865);
     data_out(1309) <= data_in(2867);
     data_out(1310) <= data_in(2873);
     data_out(1311) <= data_in(2874);
     data_out(1312) <= data_in(2875);
     data_out(1313) <= data_in(2876);
     data_out(1314) <= data_in(2878);
     data_out(1315) <= data_in(2879);
     data_out(1316) <= data_in(2881);
     data_out(1317) <= data_in(2884);
     data_out(1318) <= data_in(2885);
     data_out(1319) <= data_in(2887);
     data_out(1320) <= data_in(2889);
     data_out(1321) <= data_in(2890);
     data_out(1322) <= data_in(2892);
     data_out(1323) <= data_in(2895);
     data_out(1324) <= data_in(2897);
     data_out(1325) <= data_in(2899);
     data_out(1326) <= data_in(2907);
     data_out(1327) <= data_in(2908);
     data_out(1328) <= data_in(2910);
     data_out(1329) <= data_in(2912);
     data_out(1330) <= data_in(2913);
     data_out(1331) <= data_in(2916);
     data_out(1332) <= data_in(2917);
     data_out(1333) <= data_in(2919);
     data_out(1334) <= data_in(2921);
     data_out(1335) <= data_in(2923);
     data_out(1336) <= data_in(2924);
     data_out(1337) <= data_in(2926);
     data_out(1338) <= data_in(2927);
     data_out(1339) <= data_in(2930);
     data_out(1340) <= data_in(2931);
     data_out(1341) <= data_in(2932);
     data_out(1342) <= data_in(2933);
     data_out(1343) <= data_in(2936);
     data_out(1344) <= data_in(2937);
     data_out(1345) <= data_in(2941);
     data_out(1346) <= data_in(2945);
     data_out(1347) <= data_in(2947);
     data_out(1348) <= data_in(2948);
     data_out(1349) <= data_in(2950);
     data_out(1350) <= data_in(2954);
     data_out(1351) <= data_in(2956);
     data_out(1352) <= data_in(2959);
     data_out(1353) <= data_in(2960);
     data_out(1354) <= data_in(2964);
     data_out(1355) <= data_in(2967);
     data_out(1356) <= data_in(2970);
     data_out(1357) <= data_in(2972);
     data_out(1358) <= data_in(2973);
     data_out(1359) <= data_in(2974);
     data_out(1360) <= data_in(2975);
     data_out(1361) <= data_in(2976);
     data_out(1362) <= data_in(2981);
     data_out(1363) <= data_in(2983);
     data_out(1364) <= data_in(2988);
     data_out(1365) <= data_in(2989);
     data_out(1366) <= data_in(2991);
     data_out(1367) <= data_in(2993);
     data_out(1368) <= data_in(2995);
     data_out(1369) <= data_in(2997);
     data_out(1370) <= data_in(2998);
     data_out(1371) <= data_in(3003);
     data_out(1372) <= data_in(3006);
     data_out(1373) <= data_in(3007);
     data_out(1374) <= data_in(3011);
     data_out(1375) <= data_in(3012);
     data_out(1376) <= data_in(3015);
     data_out(1377) <= data_in(3016);
     data_out(1378) <= data_in(3020);
     data_out(1379) <= data_in(3021);
     data_out(1380) <= data_in(3022);
     data_out(1381) <= data_in(3031);
     data_out(1382) <= data_in(3033);
     data_out(1383) <= data_in(3034);
     data_out(1384) <= data_in(3037);
     data_out(1385) <= data_in(3041);
     data_out(1386) <= data_in(3044);
     data_out(1387) <= data_in(3046);
     data_out(1388) <= data_in(3050);
     data_out(1389) <= data_in(3053);
     data_out(1390) <= data_in(3054);
     data_out(1391) <= data_in(3055);
     data_out(1392) <= data_in(3061);
     data_out(1393) <= data_in(3065);
     data_out(1394) <= data_in(3066);
     data_out(1395) <= data_in(3072);
     data_out(1396) <= data_in(3073);
     data_out(1397) <= data_in(3077);
     data_out(1398) <= data_in(3081);
     data_out(1399) <= data_in(3086);
     data_out(1400) <= data_in(3088);
     data_out(1401) <= data_in(3090);
     data_out(1402) <= data_in(3095);
     data_out(1403) <= data_in(3097);
     data_out(1404) <= data_in(3100);
     data_out(1405) <= data_in(3101);
     data_out(1406) <= data_in(3107);
     data_out(1407) <= data_in(3108);
     data_out(1408) <= data_in(3115);
     data_out(1409) <= data_in(3116);
     data_out(1410) <= data_in(3126);
     data_out(1411) <= data_in(3127);
     data_out(1412) <= data_in(3128);
     data_out(1413) <= data_in(3129);
     data_out(1414) <= data_in(3133);
     data_out(1415) <= data_in(3136);
     data_out(1416) <= data_in(3138);
     data_out(1417) <= data_in(3139);
     data_out(1418) <= data_in(3140);
     data_out(1419) <= data_in(3145);
     data_out(1420) <= data_in(3147);
     data_out(1421) <= data_in(3149);
     data_out(1422) <= data_in(3150);
     data_out(1423) <= data_in(3153);
     data_out(1424) <= data_in(3154);
     data_out(1425) <= data_in(3157);
     data_out(1426) <= data_in(3162);
     data_out(1427) <= data_in(3164);
     data_out(1428) <= data_in(3165);
     data_out(1429) <= data_in(3166);
     data_out(1430) <= data_in(3170);
     data_out(1431) <= data_in(3172);
     data_out(1432) <= data_in(3174);
     data_out(1433) <= data_in(3175);
     data_out(1434) <= data_in(3179);
     data_out(1435) <= data_in(3180);
     data_out(1436) <= data_in(3181);
     data_out(1437) <= data_in(3183);
     data_out(1438) <= data_in(3184);
     data_out(1439) <= data_in(3188);
     data_out(1440) <= data_in(3191);
     data_out(1441) <= data_in(3197);
     data_out(1442) <= data_in(3198);
     data_out(1443) <= data_in(3202);
     data_out(1444) <= data_in(3203);
     data_out(1445) <= data_in(3204);
     data_out(1446) <= data_in(3205);
     data_out(1447) <= data_in(3206);
     data_out(1448) <= data_in(3208);
     data_out(1449) <= data_in(3209);
     data_out(1450) <= data_in(3210);
     data_out(1451) <= data_in(3212);
     data_out(1452) <= data_in(3213);
     data_out(1453) <= data_in(3214);
     data_out(1454) <= data_in(3215);
     data_out(1455) <= data_in(3217);
     data_out(1456) <= data_in(3218);
     data_out(1457) <= data_in(3220);
     data_out(1458) <= data_in(3222);
     data_out(1459) <= data_in(3227);
     data_out(1460) <= data_in(3228);
     data_out(1461) <= data_in(3229);
     data_out(1462) <= data_in(3232);
     data_out(1463) <= data_in(3234);
     data_out(1464) <= data_in(3235);
     data_out(1465) <= data_in(3240);
     data_out(1466) <= data_in(3247);
     data_out(1467) <= data_in(3249);
     data_out(1468) <= data_in(3251);
     data_out(1469) <= data_in(3254);
     data_out(1470) <= data_in(3255);
     data_out(1471) <= data_in(3258);
     data_out(1472) <= data_in(3259);
     data_out(1473) <= data_in(3260);
     data_out(1474) <= data_in(3264);
     data_out(1475) <= data_in(3266);
     data_out(1476) <= data_in(3267);
     data_out(1477) <= data_in(3271);
     data_out(1478) <= data_in(3274);
     data_out(1479) <= data_in(3275);
     data_out(1480) <= data_in(3277);
     data_out(1481) <= data_in(3279);
     data_out(1482) <= data_in(3282);
     data_out(1483) <= data_in(3286);
     data_out(1484) <= data_in(3287);
     data_out(1485) <= data_in(3292);
     data_out(1486) <= data_in(3293);
     data_out(1487) <= data_in(3295);
     data_out(1488) <= data_in(3297);
     data_out(1489) <= data_in(3298);
     data_out(1490) <= data_in(3300);
     data_out(1491) <= data_in(3303);
     data_out(1492) <= data_in(3304);
     data_out(1493) <= data_in(3306);
     data_out(1494) <= data_in(3307);
     data_out(1495) <= data_in(3308);
     data_out(1496) <= data_in(3309);
     data_out(1497) <= data_in(3313);
     data_out(1498) <= data_in(3314);
     data_out(1499) <= data_in(3315);
     data_out(1500) <= data_in(3316);
     data_out(1501) <= data_in(3318);
     data_out(1502) <= data_in(3321);
     data_out(1503) <= data_in(3322);
     data_out(1504) <= data_in(3324);
     data_out(1505) <= data_in(3327);
     data_out(1506) <= data_in(3328);
     data_out(1507) <= data_in(3330);
     data_out(1508) <= data_in(3331);
     data_out(1509) <= data_in(3332);
     data_out(1510) <= data_in(3338);
     data_out(1511) <= data_in(3339);
     data_out(1512) <= data_in(3342);
     data_out(1513) <= data_in(3345);
     data_out(1514) <= data_in(3349);
     data_out(1515) <= data_in(3358);
     data_out(1516) <= data_in(3359);
     data_out(1517) <= data_in(3360);
     data_out(1518) <= data_in(3361);
     data_out(1519) <= data_in(3365);
     data_out(1520) <= data_in(3372);
     data_out(1521) <= data_in(3377);
     data_out(1522) <= data_in(3383);
     data_out(1523) <= data_in(3384);
     data_out(1524) <= data_in(3393);
     data_out(1525) <= data_in(3394);
     data_out(1526) <= data_in(3397);
     data_out(1527) <= data_in(3398);
     data_out(1528) <= data_in(3402);
     data_out(1529) <= data_in(3403);
     data_out(1530) <= data_in(3409);
     data_out(1531) <= data_in(3411);
     data_out(1532) <= data_in(3412);
     data_out(1533) <= data_in(3413);
     data_out(1534) <= data_in(3414);
     data_out(1535) <= data_in(3417);
     data_out(1536) <= data_in(3419);
     data_out(1537) <= data_in(3421);
     data_out(1538) <= data_in(3425);
     data_out(1539) <= data_in(3426);
     data_out(1540) <= data_in(3427);
     data_out(1541) <= data_in(3428);
     data_out(1542) <= data_in(3429);
     data_out(1543) <= data_in(3433);
     data_out(1544) <= data_in(3435);
     data_out(1545) <= data_in(3436);
     data_out(1546) <= data_in(3437);
     data_out(1547) <= data_in(3440);
     data_out(1548) <= data_in(3448);
     data_out(1549) <= data_in(3455);
     data_out(1550) <= data_in(3456);
     data_out(1551) <= data_in(3459);
     data_out(1552) <= data_in(3466);
     data_out(1553) <= data_in(3468);
     data_out(1554) <= data_in(3472);
     data_out(1555) <= data_in(3474);
     data_out(1556) <= data_in(3475);
     data_out(1557) <= data_in(3477);
     data_out(1558) <= data_in(3478);
     data_out(1559) <= data_in(3479);
     data_out(1560) <= data_in(3484);
     data_out(1561) <= data_in(3488);
     data_out(1562) <= data_in(3491);
     data_out(1563) <= data_in(3492);
     data_out(1564) <= data_in(3494);
     data_out(1565) <= data_in(3495);
     data_out(1566) <= data_in(3497);
     data_out(1567) <= data_in(3498);
     data_out(1568) <= data_in(3504);
     data_out(1569) <= data_in(3508);
     data_out(1570) <= data_in(3510);
     data_out(1571) <= data_in(3513);
     data_out(1572) <= data_in(3517);
     data_out(1573) <= data_in(3521);
     data_out(1574) <= data_in(3523);
     data_out(1575) <= data_in(3525);
     data_out(1576) <= data_in(3528);
     data_out(1577) <= data_in(3530);
     data_out(1578) <= data_in(3532);
     data_out(1579) <= data_in(3533);
     data_out(1580) <= data_in(3538);
     data_out(1581) <= data_in(3550);
     data_out(1582) <= data_in(3551);
     data_out(1583) <= data_in(3553);
     data_out(1584) <= data_in(3560);
     data_out(1585) <= data_in(3561);
     data_out(1586) <= data_in(3564);
     data_out(1587) <= data_in(3568);
     data_out(1588) <= data_in(3570);
     data_out(1589) <= data_in(3571);
     data_out(1590) <= data_in(3574);
     data_out(1591) <= data_in(3575);
     data_out(1592) <= data_in(3576);
     data_out(1593) <= data_in(3585);
     data_out(1594) <= data_in(3587);
     data_out(1595) <= data_in(3588);
     data_out(1596) <= data_in(3589);
     data_out(1597) <= data_in(3590);
     data_out(1598) <= data_in(3591);
     data_out(1599) <= data_in(3592);
     data_out(1600) <= data_in(3596);
     data_out(1601) <= data_in(3597);
     data_out(1602) <= data_in(3600);
     data_out(1603) <= data_in(3606);
     data_out(1604) <= data_in(3607);
     data_out(1605) <= data_in(3608);
     data_out(1606) <= data_in(3613);
     data_out(1607) <= data_in(3615);
     data_out(1608) <= data_in(3617);
     data_out(1609) <= data_in(3622);
     data_out(1610) <= data_in(3624);
     data_out(1611) <= data_in(3629);
     data_out(1612) <= data_in(3631);
     data_out(1613) <= data_in(3632);
     data_out(1614) <= data_in(3634);
     data_out(1615) <= data_in(3635);
     data_out(1616) <= data_in(3638);
     data_out(1617) <= data_in(3639);
     data_out(1618) <= data_in(3640);
     data_out(1619) <= data_in(3648);
     data_out(1620) <= data_in(3649);
     data_out(1621) <= data_in(3651);
     data_out(1622) <= data_in(3657);
     data_out(1623) <= data_in(3660);
     data_out(1624) <= data_in(3661);
     data_out(1625) <= data_in(3664);
     data_out(1626) <= data_in(3670);
     data_out(1627) <= data_in(3671);
     data_out(1628) <= data_in(3672);
     data_out(1629) <= data_in(3674);
     data_out(1630) <= data_in(3676);
     data_out(1631) <= data_in(3677);
     data_out(1632) <= data_in(3678);
     data_out(1633) <= data_in(3684);
     data_out(1634) <= data_in(3686);
     data_out(1635) <= data_in(3692);
     data_out(1636) <= data_in(3694);
     data_out(1637) <= data_in(3695);
     data_out(1638) <= data_in(3697);
     data_out(1639) <= data_in(3699);
     data_out(1640) <= data_in(3700);
     data_out(1641) <= data_in(3701);
     data_out(1642) <= data_in(3702);
     data_out(1643) <= data_in(3706);
     data_out(1644) <= data_in(3707);
     data_out(1645) <= data_in(3708);
     data_out(1646) <= data_in(3710);
     data_out(1647) <= data_in(3712);
     data_out(1648) <= data_in(3714);
     data_out(1649) <= data_in(3717);
     data_out(1650) <= data_in(3718);
     data_out(1651) <= data_in(3723);
     data_out(1652) <= data_in(3724);
     data_out(1653) <= data_in(3725);
     data_out(1654) <= data_in(3732);
     data_out(1655) <= data_in(3734);
     data_out(1656) <= data_in(3737);
     data_out(1657) <= data_in(3739);
     data_out(1658) <= data_in(3740);
     data_out(1659) <= data_in(3742);
     data_out(1660) <= data_in(3744);
     data_out(1661) <= data_in(3746);
     data_out(1662) <= data_in(3750);
     data_out(1663) <= data_in(3751);
     data_out(1664) <= data_in(3755);
     data_out(1665) <= data_in(3756);
     data_out(1666) <= data_in(3759);
     data_out(1667) <= data_in(3761);
     data_out(1668) <= data_in(3765);
     data_out(1669) <= data_in(3768);
     data_out(1670) <= data_in(3772);
     data_out(1671) <= data_in(3775);
     data_out(1672) <= data_in(3776);
     data_out(1673) <= data_in(3781);
     data_out(1674) <= data_in(3782);
     data_out(1675) <= data_in(3783);
     data_out(1676) <= data_in(3789);
     data_out(1677) <= data_in(3790);
     data_out(1678) <= data_in(3793);
     data_out(1679) <= data_in(3794);
     data_out(1680) <= data_in(3798);
     data_out(1681) <= data_in(3801);
     data_out(1682) <= data_in(3803);
     data_out(1683) <= data_in(3805);
     data_out(1684) <= data_in(3806);
     data_out(1685) <= data_in(3808);
     data_out(1686) <= data_in(3809);
     data_out(1687) <= data_in(3810);
     data_out(1688) <= data_in(3819);
     data_out(1689) <= data_in(3821);
     data_out(1690) <= data_in(3824);
     data_out(1691) <= data_in(3829);
     data_out(1692) <= data_in(3831);
     data_out(1693) <= data_in(3839);
     data_out(1694) <= data_in(3842);
     data_out(1695) <= data_in(3844);
     data_out(1696) <= data_in(3845);
     data_out(1697) <= data_in(3848);
     data_out(1698) <= data_in(3850);
     data_out(1699) <= data_in(3851);
     data_out(1700) <= data_in(3852);
     data_out(1701) <= data_in(3855);
     data_out(1702) <= data_in(3856);
     data_out(1703) <= data_in(3858);
     data_out(1704) <= data_in(3860);
     data_out(1705) <= data_in(3861);
     data_out(1706) <= data_in(3862);
     data_out(1707) <= data_in(3863);
     data_out(1708) <= data_in(3864);
     data_out(1709) <= data_in(3868);
     data_out(1710) <= data_in(3869);
     data_out(1711) <= data_in(3874);
     data_out(1712) <= data_in(3877);
     data_out(1713) <= data_in(3879);
     data_out(1714) <= data_in(3883);
     data_out(1715) <= data_in(3884);
     data_out(1716) <= data_in(3888);
     data_out(1717) <= data_in(3889);
     data_out(1718) <= data_in(3891);
     data_out(1719) <= data_in(3894);
     data_out(1720) <= data_in(3895);
     data_out(1721) <= data_in(3897);
     data_out(1722) <= data_in(3902);
     data_out(1723) <= data_in(3903);
     data_out(1724) <= data_in(3906);
     data_out(1725) <= data_in(3910);
     data_out(1726) <= data_in(3911);
     data_out(1727) <= data_in(3922);
     data_out(1728) <= data_in(3923);
     data_out(1729) <= data_in(3927);
     data_out(1730) <= data_in(3930);
     data_out(1731) <= data_in(3931);
     data_out(1732) <= data_in(3932);
     data_out(1733) <= data_in(3934);
     data_out(1734) <= data_in(3935);
     data_out(1735) <= data_in(3939);
     data_out(1736) <= data_in(3941);
     data_out(1737) <= data_in(3942);
     data_out(1738) <= data_in(3943);
     data_out(1739) <= data_in(3945);
     data_out(1740) <= data_in(3951);
     data_out(1741) <= data_in(3952);
     data_out(1742) <= data_in(3953);
     data_out(1743) <= data_in(3956);
     data_out(1744) <= data_in(3958);
     data_out(1745) <= data_in(3961);
     data_out(1746) <= data_in(3962);
     data_out(1747) <= data_in(3964);
     data_out(1748) <= data_in(3966);
     data_out(1749) <= data_in(3967);
     data_out(1750) <= data_in(3969);
     data_out(1751) <= data_in(3973);
     data_out(1752) <= data_in(3976);
     data_out(1753) <= data_in(3978);
     data_out(1754) <= data_in(3979);
     data_out(1755) <= data_in(3981);
     data_out(1756) <= data_in(3984);
     data_out(1757) <= data_in(3985);
     data_out(1758) <= data_in(3990);
     data_out(1759) <= data_in(3991);
     data_out(1760) <= data_in(3993);
     data_out(1761) <= data_in(3996);
     data_out(1762) <= data_in(4000);
     data_out(1763) <= data_in(4003);
     data_out(1764) <= data_in(4004);
     data_out(1765) <= data_in(4005);
     data_out(1766) <= data_in(4006);
     data_out(1767) <= data_in(4010);
     data_out(1768) <= data_in(4012);
     data_out(1769) <= data_in(4014);
     data_out(1770) <= data_in(4022);
     data_out(1771) <= data_in(4024);
     data_out(1772) <= data_in(4028);
     data_out(1773) <= data_in(4029);
     data_out(1774) <= data_in(4035);
     data_out(1775) <= data_in(4037);
     data_out(1776) <= data_in(4042);
     data_out(1777) <= data_in(4046);
     data_out(1778) <= data_in(4047);
     data_out(1779) <= data_in(4056);
     data_out(1780) <= data_in(4061);
     data_out(1781) <= data_in(4065);
     data_out(1782) <= data_in(4070);
     data_out(1783) <= data_in(4071);
     data_out(1784) <= data_in(4073);
     data_out(1785) <= data_in(4074);
     data_out(1786) <= data_in(4078);
     data_out(1787) <= data_in(4081);
     data_out(1788) <= data_in(4089);
     data_out(1789) <= data_in(4094);
     data_out(1790) <= data_in(4096);
     data_out(1791) <= data_in(4097);
     data_out(1792) <= data_in(4098);
     data_out(1793) <= data_in(4099);
     data_out(1794) <= data_in(4103);
     data_out(1795) <= data_in(4106);
     data_out(1796) <= data_in(4110);
     data_out(1797) <= data_in(4111);
     data_out(1798) <= data_in(4112);
     data_out(1799) <= data_in(4113);
     data_out(1800) <= data_in(4116);
     data_out(1801) <= data_in(4118);
     data_out(1802) <= data_in(4119);
     data_out(1803) <= data_in(4122);
     data_out(1804) <= data_in(4124);
     data_out(1805) <= data_in(4125);
     data_out(1806) <= data_in(4126);
     data_out(1807) <= data_in(4129);
     data_out(1808) <= data_in(4130);
     data_out(1809) <= data_in(4131);
     data_out(1810) <= data_in(4134);
     data_out(1811) <= data_in(4135);
     data_out(1812) <= data_in(4136);
     data_out(1813) <= data_in(4139);
     data_out(1814) <= data_in(4140);
     data_out(1815) <= data_in(4141);
     data_out(1816) <= data_in(4142);
     data_out(1817) <= data_in(4146);
     data_out(1818) <= data_in(4148);
     data_out(1819) <= data_in(4159);
     data_out(1820) <= data_in(4161);
     data_out(1821) <= data_in(4165);
     data_out(1822) <= data_in(4166);
     data_out(1823) <= data_in(4171);
     data_out(1824) <= data_in(4173);
     data_out(1825) <= data_in(4174);
     data_out(1826) <= data_in(4181);
     data_out(1827) <= data_in(4182);
     data_out(1828) <= data_in(4184);
     data_out(1829) <= data_in(4185);
     data_out(1830) <= data_in(4186);
     data_out(1831) <= data_in(4188);
     data_out(1832) <= data_in(4190);
     data_out(1833) <= data_in(4193);
     data_out(1834) <= data_in(4204);
     data_out(1835) <= data_in(4207);
     data_out(1836) <= data_in(4210);
     data_out(1837) <= data_in(4212);
     data_out(1838) <= data_in(4216);
     data_out(1839) <= data_in(4219);
     data_out(1840) <= data_in(4220);
     data_out(1841) <= data_in(4223);
     data_out(1842) <= data_in(4224);
     data_out(1843) <= data_in(4230);
     data_out(1844) <= data_in(4232);
     data_out(1845) <= data_in(4233);
     data_out(1846) <= data_in(4234);
     data_out(1847) <= data_in(4236);
     data_out(1848) <= data_in(4237);
     data_out(1849) <= data_in(4240);
     data_out(1850) <= data_in(4241);
     data_out(1851) <= data_in(4244);
     data_out(1852) <= data_in(4245);
     data_out(1853) <= data_in(4246);
     data_out(1854) <= data_in(4249);
     data_out(1855) <= data_in(4251);
     data_out(1856) <= data_in(4252);
     data_out(1857) <= data_in(4254);
     data_out(1858) <= data_in(4260);
     data_out(1859) <= data_in(4267);
     data_out(1860) <= data_in(4270);
     data_out(1861) <= data_in(4271);
     data_out(1862) <= data_in(4274);
     data_out(1863) <= data_in(4276);
     data_out(1864) <= data_in(4277);
     data_out(1865) <= data_in(4279);
     data_out(1866) <= data_in(4282);
     data_out(1867) <= data_in(4283);
     data_out(1868) <= data_in(4284);
     data_out(1869) <= data_in(4288);
     data_out(1870) <= data_in(4289);
     data_out(1871) <= data_in(4294);
     data_out(1872) <= data_in(4297);
     data_out(1873) <= data_in(4298);
     data_out(1874) <= data_in(4302);
     data_out(1875) <= data_in(4304);
     data_out(1876) <= data_in(4305);
     data_out(1877) <= data_in(4306);
     data_out(1878) <= data_in(4309);
     data_out(1879) <= data_in(4317);
     data_out(1880) <= data_in(4329);
     data_out(1881) <= data_in(4330);
     data_out(1882) <= data_in(4332);
     data_out(1883) <= data_in(4337);
     data_out(1884) <= data_in(4339);
     data_out(1885) <= data_in(4340);
     data_out(1886) <= data_in(4342);
     data_out(1887) <= data_in(4345);
     data_out(1888) <= data_in(4346);
     data_out(1889) <= data_in(4350);
     data_out(1890) <= data_in(4354);
     data_out(1891) <= data_in(4358);
     data_out(1892) <= data_in(4359);
     data_out(1893) <= data_in(4360);
     data_out(1894) <= data_in(4363);
     data_out(1895) <= data_in(4368);
     data_out(1896) <= data_in(4369);
     data_out(1897) <= data_in(4372);
     data_out(1898) <= data_in(4375);
     data_out(1899) <= data_in(4377);
     data_out(1900) <= data_in(4379);
     data_out(1901) <= data_in(4380);
     data_out(1902) <= data_in(4383);
     data_out(1903) <= data_in(4384);
     data_out(1904) <= data_in(4385);
     data_out(1905) <= data_in(4391);
     data_out(1906) <= data_in(4402);
     data_out(1907) <= data_in(4406);
     data_out(1908) <= data_in(4412);
     data_out(1909) <= data_in(4416);
     data_out(1910) <= data_in(4417);
     data_out(1911) <= data_in(4418);
     data_out(1912) <= data_in(4420);
     data_out(1913) <= data_in(4422);
     data_out(1914) <= data_in(4425);
     data_out(1915) <= data_in(4426);
     data_out(1916) <= data_in(4429);
     data_out(1917) <= data_in(4435);
     data_out(1918) <= data_in(4439);
     data_out(1919) <= data_in(4442);
     data_out(1920) <= data_in(4446);
     data_out(1921) <= data_in(4447);
     data_out(1922) <= data_in(4448);
     data_out(1923) <= data_in(4453);
     data_out(1924) <= data_in(4454);
     data_out(1925) <= data_in(4456);
     data_out(1926) <= data_in(4457);
     data_out(1927) <= data_in(4458);
     data_out(1928) <= data_in(4459);
     data_out(1929) <= data_in(4461);
     data_out(1930) <= data_in(4467);
     data_out(1931) <= data_in(4468);
     data_out(1932) <= data_in(4473);
     data_out(1933) <= data_in(4474);
     data_out(1934) <= data_in(4475);
     data_out(1935) <= data_in(4478);
     data_out(1936) <= data_in(4479);
     data_out(1937) <= data_in(4480);
     data_out(1938) <= data_in(4483);
     data_out(1939) <= data_in(4484);
     data_out(1940) <= data_in(4485);
     data_out(1941) <= data_in(4495);
     data_out(1942) <= data_in(4496);
     data_out(1943) <= data_in(4497);
     data_out(1944) <= data_in(4499);
     data_out(1945) <= data_in(4500);
     data_out(1946) <= data_in(4501);
     data_out(1947) <= data_in(4503);
     data_out(1948) <= data_in(4505);
     data_out(1949) <= data_in(4508);
     data_out(1950) <= data_in(4510);
     data_out(1951) <= data_in(4513);
     data_out(1952) <= data_in(4516);
     data_out(1953) <= data_in(4518);
     data_out(1954) <= data_in(4522);
     data_out(1955) <= data_in(4524);
     data_out(1956) <= data_in(4528);
     data_out(1957) <= data_in(4529);
     data_out(1958) <= data_in(4532);
     data_out(1959) <= data_in(4534);
     data_out(1960) <= data_in(4535);
     data_out(1961) <= data_in(4538);
     data_out(1962) <= data_in(4539);
     data_out(1963) <= data_in(4541);
     data_out(1964) <= data_in(4543);
     data_out(1965) <= data_in(4545);
     data_out(1966) <= data_in(4551);
     data_out(1967) <= data_in(4554);
     data_out(1968) <= data_in(4558);
     data_out(1969) <= data_in(4560);
     data_out(1970) <= data_in(4564);
     data_out(1971) <= data_in(4565);
     data_out(1972) <= data_in(4567);
     data_out(1973) <= data_in(4568);
     data_out(1974) <= data_in(4569);
     data_out(1975) <= data_in(4570);
     data_out(1976) <= data_in(4571);
     data_out(1977) <= data_in(4573);
     data_out(1978) <= data_in(4575);
     data_out(1979) <= data_in(4576);
     data_out(1980) <= data_in(4579);
     data_out(1981) <= data_in(4582);
     data_out(1982) <= data_in(4584);
     data_out(1983) <= data_in(4586);
     data_out(1984) <= data_in(4589);
     data_out(1985) <= data_in(4594);
     data_out(1986) <= data_in(4596);
     data_out(1987) <= data_in(4599);
     data_out(1988) <= data_in(4607);
     data_out(1989) <= data_in(4608);
     data_out(1990) <= data_in(4609);
     data_out(1991) <= data_in(4612);
     data_out(1992) <= data_in(4613);
     data_out(1993) <= data_in(4616);
     data_out(1994) <= data_in(4622);
     data_out(1995) <= data_in(4623);
     data_out(1996) <= data_in(4624);
     data_out(1997) <= data_in(4625);
     data_out(1998) <= data_in(4626);
     data_out(1999) <= data_in(4628);
     data_out(2000) <= data_in(4635);
     data_out(2001) <= data_in(4637);
     data_out(2002) <= data_in(4638);
     data_out(2003) <= data_in(4641);
     data_out(2004) <= data_in(4644);
     data_out(2005) <= data_in(4645);
     data_out(2006) <= data_in(4646);
     data_out(2007) <= data_in(4649);
     data_out(2008) <= data_in(4651);
     data_out(2009) <= data_in(4653);
     data_out(2010) <= data_in(4654);
     data_out(2011) <= data_in(4656);
     data_out(2012) <= data_in(4657);
     data_out(2013) <= data_in(4659);
     data_out(2014) <= data_in(4660);
     data_out(2015) <= data_in(4663);
     data_out(2016) <= data_in(4665);
     data_out(2017) <= data_in(4672);
     data_out(2018) <= data_in(4674);
     data_out(2019) <= data_in(4675);
     data_out(2020) <= data_in(4677);
     data_out(2021) <= data_in(4686);
     data_out(2022) <= data_in(4689);
     data_out(2023) <= data_in(4694);
     data_out(2024) <= data_in(4696);
     data_out(2025) <= data_in(4697);
     data_out(2026) <= data_in(4698);
     data_out(2027) <= data_in(4702);
     data_out(2028) <= data_in(4704);
     data_out(2029) <= data_in(4705);
     data_out(2030) <= data_in(4710);
     data_out(2031) <= data_in(4711);
     data_out(2032) <= data_in(4712);
     data_out(2033) <= data_in(4713);
     data_out(2034) <= data_in(4715);
     data_out(2035) <= data_in(4716);
     data_out(2036) <= data_in(4718);
     data_out(2037) <= data_in(4719);
     data_out(2038) <= data_in(4720);
     data_out(2039) <= data_in(4723);
     data_out(2040) <= data_in(4724);
     data_out(2041) <= data_in(4725);
     data_out(2042) <= data_in(4726);
     data_out(2043) <= data_in(4731);
     data_out(2044) <= data_in(4732);
     data_out(2045) <= data_in(4739);
     data_out(2046) <= data_in(4741);
     data_out(2047) <= data_in(4744);
     data_out(2048) <= data_in(4745);
     data_out(2049) <= data_in(4746);
     data_out(2050) <= data_in(4747);
     data_out(2051) <= data_in(4750);
     data_out(2052) <= data_in(4751);
     data_out(2053) <= data_in(4754);
     data_out(2054) <= data_in(4755);
     data_out(2055) <= data_in(4756);
     data_out(2056) <= data_in(4758);
     data_out(2057) <= data_in(4760);
     data_out(2058) <= data_in(4761);
     data_out(2059) <= data_in(4763);
     data_out(2060) <= data_in(4765);
     data_out(2061) <= data_in(4768);
     data_out(2062) <= data_in(4769);
     data_out(2063) <= data_in(4771);
     data_out(2064) <= data_in(4773);
     data_out(2065) <= data_in(4775);
     data_out(2066) <= data_in(4777);
     data_out(2067) <= data_in(4780);
     data_out(2068) <= data_in(4782);
     data_out(2069) <= data_in(4783);
     data_out(2070) <= data_in(4785);
     data_out(2071) <= data_in(4793);
     data_out(2072) <= data_in(4794);
     data_out(2073) <= data_in(4801);
     data_out(2074) <= data_in(4804);
     data_out(2075) <= data_in(4809);
     data_out(2076) <= data_in(4810);
     data_out(2077) <= data_in(4812);
     data_out(2078) <= data_in(4817);
     data_out(2079) <= data_in(4820);
     data_out(2080) <= data_in(4822);
     data_out(2081) <= data_in(4823);
     data_out(2082) <= data_in(4826);
     data_out(2083) <= data_in(4827);
     data_out(2084) <= data_in(4829);
     data_out(2085) <= data_in(4835);
     data_out(2086) <= data_in(4842);
     data_out(2087) <= data_in(4844);
     data_out(2088) <= data_in(4845);
     data_out(2089) <= data_in(4846);
     data_out(2090) <= data_in(4857);
     data_out(2091) <= data_in(4859);
     data_out(2092) <= data_in(4862);
     data_out(2093) <= data_in(4864);
     data_out(2094) <= data_in(4865);
     data_out(2095) <= data_in(4866);
     data_out(2096) <= data_in(4867);
     data_out(2097) <= data_in(4871);
     data_out(2098) <= data_in(4875);
     data_out(2099) <= data_in(4879);
     data_out(2100) <= data_in(4883);
     data_out(2101) <= data_in(4887);
     data_out(2102) <= data_in(4890);
     data_out(2103) <= data_in(4891);
     data_out(2104) <= data_in(4892);
     data_out(2105) <= data_in(4893);
     data_out(2106) <= data_in(4895);
     data_out(2107) <= data_in(4896);
     data_out(2108) <= data_in(4900);
     data_out(2109) <= data_in(4901);
     data_out(2110) <= data_in(4902);
     data_out(2111) <= data_in(4904);
     data_out(2112) <= data_in(4907);
     data_out(2113) <= data_in(4909);
     data_out(2114) <= data_in(4911);
     data_out(2115) <= data_in(4915);
     data_out(2116) <= data_in(4916);
     data_out(2117) <= data_in(4918);
     data_out(2118) <= data_in(4921);
     data_out(2119) <= data_in(4922);
     data_out(2120) <= data_in(4923);
     data_out(2121) <= data_in(4924);
     data_out(2122) <= data_in(4927);
     data_out(2123) <= data_in(4931);
     data_out(2124) <= data_in(4932);
     data_out(2125) <= data_in(4933);
     data_out(2126) <= data_in(4934);
     data_out(2127) <= data_in(4938);
     data_out(2128) <= data_in(4939);
     data_out(2129) <= data_in(4941);
     data_out(2130) <= data_in(4944);
     data_out(2131) <= data_in(4945);
     data_out(2132) <= data_in(4946);
     data_out(2133) <= data_in(4947);
     data_out(2134) <= data_in(4949);
     data_out(2135) <= data_in(4953);
     data_out(2136) <= data_in(4956);
     data_out(2137) <= data_in(4958);
     data_out(2138) <= data_in(4959);
     data_out(2139) <= data_in(4962);
     data_out(2140) <= data_in(4968);
     data_out(2141) <= data_in(4970);
     data_out(2142) <= data_in(4975);
     data_out(2143) <= data_in(4976);
     data_out(2144) <= data_in(4977);
     data_out(2145) <= data_in(4983);
     data_out(2146) <= data_in(4987);
     data_out(2147) <= data_in(4988);
     data_out(2148) <= data_in(4990);
     data_out(2149) <= data_in(4993);
     data_out(2150) <= data_in(4999);
     data_out(2151) <= data_in(5001);
     data_out(2152) <= data_in(5007);
     data_out(2153) <= data_in(5013);
     data_out(2154) <= data_in(5014);
     data_out(2155) <= data_in(5015);
     data_out(2156) <= data_in(5020);
     data_out(2157) <= data_in(5023);
     data_out(2158) <= data_in(5027);
     data_out(2159) <= data_in(5028);
     data_out(2160) <= data_in(5030);
     data_out(2161) <= data_in(5031);
     data_out(2162) <= data_in(5033);
     data_out(2163) <= data_in(5034);
     data_out(2164) <= data_in(5035);
     data_out(2165) <= data_in(5040);
     data_out(2166) <= data_in(5041);
     data_out(2167) <= data_in(5042);
     data_out(2168) <= data_in(5046);
     data_out(2169) <= data_in(5049);
     data_out(2170) <= data_in(5050);
     data_out(2171) <= data_in(5051);
     data_out(2172) <= data_in(5052);
     data_out(2173) <= data_in(5054);
     data_out(2174) <= data_in(5062);
     data_out(2175) <= data_in(5066);
     data_out(2176) <= data_in(5067);
     data_out(2177) <= data_in(5069);
     data_out(2178) <= data_in(5072);
     data_out(2179) <= data_in(5082);
     data_out(2180) <= data_in(5087);
     data_out(2181) <= data_in(5089);
     data_out(2182) <= data_in(5090);
     data_out(2183) <= data_in(5091);
     data_out(2184) <= data_in(5093);
     data_out(2185) <= data_in(5097);
     data_out(2186) <= data_in(5098);
     data_out(2187) <= data_in(5100);
     data_out(2188) <= data_in(5104);
     data_out(2189) <= data_in(5109);
     data_out(2190) <= data_in(5110);
     data_out(2191) <= data_in(5111);
     data_out(2192) <= data_in(5114);
     data_out(2193) <= data_in(5116);
     data_out(2194) <= data_in(5117);
     data_out(2195) <= data_in(5118);
     data_out(2196) <= data_in(5123);
     data_out(2197) <= data_in(5131);
     data_out(2198) <= data_in(5133);
     data_out(2199) <= data_in(5135);
     data_out(2200) <= data_in(5141);
     data_out(2201) <= data_in(5143);
     data_out(2202) <= data_in(5144);
     data_out(2203) <= data_in(5145);
     data_out(2204) <= data_in(5146);
     data_out(2205) <= data_in(5149);
     data_out(2206) <= data_in(5151);
     data_out(2207) <= data_in(5152);
     data_out(2208) <= data_in(5154);
     data_out(2209) <= data_in(5155);
     data_out(2210) <= data_in(5157);
     data_out(2211) <= data_in(5158);
     data_out(2212) <= data_in(5159);
     data_out(2213) <= data_in(5160);
     data_out(2214) <= data_in(5168);
     data_out(2215) <= data_in(5169);
     data_out(2216) <= data_in(5171);
     data_out(2217) <= data_in(5174);
     data_out(2218) <= data_in(5176);
     data_out(2219) <= data_in(5179);
     data_out(2220) <= data_in(5180);
     data_out(2221) <= data_in(5181);
     data_out(2222) <= data_in(5182);
     data_out(2223) <= data_in(5184);
     data_out(2224) <= data_in(5187);
     data_out(2225) <= data_in(5190);
     data_out(2226) <= data_in(5195);
     data_out(2227) <= data_in(5196);
     data_out(2228) <= data_in(5199);
     data_out(2229) <= data_in(5201);
     data_out(2230) <= data_in(5205);
     data_out(2231) <= data_in(5206);
     data_out(2232) <= data_in(5207);
     data_out(2233) <= data_in(5211);
     data_out(2234) <= data_in(5214);
     data_out(2235) <= data_in(5216);
     data_out(2236) <= data_in(5219);
     data_out(2237) <= data_in(5226);
     data_out(2238) <= data_in(5227);
     data_out(2239) <= data_in(5228);
     data_out(2240) <= data_in(5230);
     data_out(2241) <= data_in(5233);
     data_out(2242) <= data_in(5234);
     data_out(2243) <= data_in(5235);
     data_out(2244) <= data_in(5236);
     data_out(2245) <= data_in(5237);
     data_out(2246) <= data_in(5240);
     data_out(2247) <= data_in(5243);
     data_out(2248) <= data_in(5244);
     data_out(2249) <= data_in(5246);
     data_out(2250) <= data_in(5249);
     data_out(2251) <= data_in(5251);
     data_out(2252) <= data_in(5252);
     data_out(2253) <= data_in(5253);
     data_out(2254) <= data_in(5255);
     data_out(2255) <= data_in(5256);
     data_out(2256) <= data_in(5260);
     data_out(2257) <= data_in(5263);
     data_out(2258) <= data_in(5265);
     data_out(2259) <= data_in(5267);
     data_out(2260) <= data_in(5268);
     data_out(2261) <= data_in(5269);
     data_out(2262) <= data_in(5271);
     data_out(2263) <= data_in(5280);
     data_out(2264) <= data_in(5281);
     data_out(2265) <= data_in(5284);
     data_out(2266) <= data_in(5286);
     data_out(2267) <= data_in(5287);
     data_out(2268) <= data_in(5288);
     data_out(2269) <= data_in(5290);
     data_out(2270) <= data_in(5291);
     data_out(2271) <= data_in(5298);
     data_out(2272) <= data_in(5305);
     data_out(2273) <= data_in(5309);
     data_out(2274) <= data_in(5314);
     data_out(2275) <= data_in(5315);
     data_out(2276) <= data_in(5318);
     data_out(2277) <= data_in(5320);
     data_out(2278) <= data_in(5321);
     data_out(2279) <= data_in(5326);
     data_out(2280) <= data_in(5327);
     data_out(2281) <= data_in(5328);
     data_out(2282) <= data_in(5331);
     data_out(2283) <= data_in(5336);
     data_out(2284) <= data_in(5339);
     data_out(2285) <= data_in(5340);
     data_out(2286) <= data_in(5343);
     data_out(2287) <= data_in(5347);
     data_out(2288) <= data_in(5348);
     data_out(2289) <= data_in(5349);
     data_out(2290) <= data_in(5356);
     data_out(2291) <= data_in(5357);
     data_out(2292) <= data_in(5359);
     data_out(2293) <= data_in(5361);
     data_out(2294) <= data_in(5363);
     data_out(2295) <= data_in(5367);
     data_out(2296) <= data_in(5373);
     data_out(2297) <= data_in(5374);
     data_out(2298) <= data_in(5375);
     data_out(2299) <= data_in(5380);
     data_out(2300) <= data_in(5381);
     data_out(2301) <= data_in(5382);
     data_out(2302) <= data_in(5384);
     data_out(2303) <= data_in(5385);
     data_out(2304) <= data_in(5387);
     data_out(2305) <= data_in(5390);
     data_out(2306) <= data_in(5395);
     data_out(2307) <= data_in(5399);
     data_out(2308) <= data_in(5400);
     data_out(2309) <= data_in(5401);
     data_out(2310) <= data_in(5403);
     data_out(2311) <= data_in(5404);
     data_out(2312) <= data_in(5406);
     data_out(2313) <= data_in(5411);
     data_out(2314) <= data_in(5415);
     data_out(2315) <= data_in(5416);
     data_out(2316) <= data_in(5419);
     data_out(2317) <= data_in(5420);
     data_out(2318) <= data_in(5421);
     data_out(2319) <= data_in(5423);
     data_out(2320) <= data_in(5425);
     data_out(2321) <= data_in(5426);
     data_out(2322) <= data_in(5427);
     data_out(2323) <= data_in(5428);
     data_out(2324) <= data_in(5429);
     data_out(2325) <= data_in(5433);
     data_out(2326) <= data_in(5435);
     data_out(2327) <= data_in(5437);
     data_out(2328) <= data_in(5442);
     data_out(2329) <= data_in(5443);
     data_out(2330) <= data_in(5446);
     data_out(2331) <= data_in(5453);
     data_out(2332) <= data_in(5458);
     data_out(2333) <= data_in(5460);
     data_out(2334) <= data_in(5461);
     data_out(2335) <= data_in(5462);
     data_out(2336) <= data_in(5463);
     data_out(2337) <= data_in(5470);
     data_out(2338) <= data_in(5471);
     data_out(2339) <= data_in(5474);
     data_out(2340) <= data_in(5475);
     data_out(2341) <= data_in(5476);
     data_out(2342) <= data_in(5477);
     data_out(2343) <= data_in(5478);
     data_out(2344) <= data_in(5482);
     data_out(2345) <= data_in(5484);
     data_out(2346) <= data_in(5487);
     data_out(2347) <= data_in(5488);
     data_out(2348) <= data_in(5489);
     data_out(2349) <= data_in(5496);
     data_out(2350) <= data_in(5497);
     data_out(2351) <= data_in(5498);
     data_out(2352) <= data_in(5501);
     data_out(2353) <= data_in(5502);
     data_out(2354) <= data_in(5503);
     data_out(2355) <= data_in(5505);
     data_out(2356) <= data_in(5506);
     data_out(2357) <= data_in(5508);
     data_out(2358) <= data_in(5510);
     data_out(2359) <= data_in(5511);
     data_out(2360) <= data_in(5513);
     data_out(2361) <= data_in(5514);
     data_out(2362) <= data_in(5519);
     data_out(2363) <= data_in(5520);
     data_out(2364) <= data_in(5524);
     data_out(2365) <= data_in(5525);
     data_out(2366) <= data_in(5528);
     data_out(2367) <= data_in(5529);
     data_out(2368) <= data_in(5530);
     data_out(2369) <= data_in(5532);
     data_out(2370) <= data_in(5534);
     data_out(2371) <= data_in(5535);
     data_out(2372) <= data_in(5540);
     data_out(2373) <= data_in(5541);
     data_out(2374) <= data_in(5542);
     data_out(2375) <= data_in(5544);
     data_out(2376) <= data_in(5547);
     data_out(2377) <= data_in(5548);
     data_out(2378) <= data_in(5551);
     data_out(2379) <= data_in(5554);
     data_out(2380) <= data_in(5555);
     data_out(2381) <= data_in(5556);
     data_out(2382) <= data_in(5558);
     data_out(2383) <= data_in(5560);
     data_out(2384) <= data_in(5563);
     data_out(2385) <= data_in(5564);
     data_out(2386) <= data_in(5566);
     data_out(2387) <= data_in(5567);
     data_out(2388) <= data_in(5568);
     data_out(2389) <= data_in(5570);
     data_out(2390) <= data_in(5571);
     data_out(2391) <= data_in(5574);
     data_out(2392) <= data_in(5581);
     data_out(2393) <= data_in(5582);
     data_out(2394) <= data_in(5583);
     data_out(2395) <= data_in(5585);
     data_out(2396) <= data_in(5586);
     data_out(2397) <= data_in(5588);
     data_out(2398) <= data_in(5590);
     data_out(2399) <= data_in(5591);
     data_out(2400) <= data_in(5592);
     data_out(2401) <= data_in(5594);
     data_out(2402) <= data_in(5595);
     data_out(2403) <= data_in(5596);
     data_out(2404) <= data_in(5597);
     data_out(2405) <= data_in(5600);
     data_out(2406) <= data_in(5605);
     data_out(2407) <= data_in(5607);
     data_out(2408) <= data_in(5610);
     data_out(2409) <= data_in(5613);
     data_out(2410) <= data_in(5616);
     data_out(2411) <= data_in(5619);
     data_out(2412) <= data_in(5621);
     data_out(2413) <= data_in(5625);
     data_out(2414) <= data_in(5627);
     data_out(2415) <= data_in(5634);
     data_out(2416) <= data_in(5635);
     data_out(2417) <= data_in(5637);
     data_out(2418) <= data_in(5638);
     data_out(2419) <= data_in(5639);
     data_out(2420) <= data_in(5641);
     data_out(2421) <= data_in(5642);
     data_out(2422) <= data_in(5643);
     data_out(2423) <= data_in(5644);
     data_out(2424) <= data_in(5646);
     data_out(2425) <= data_in(5648);
     data_out(2426) <= data_in(5649);
     data_out(2427) <= data_in(5651);
     data_out(2428) <= data_in(5653);
     data_out(2429) <= data_in(5654);
     data_out(2430) <= data_in(5655);
     data_out(2431) <= data_in(5658);
     data_out(2432) <= data_in(5662);
     data_out(2433) <= data_in(5665);
     data_out(2434) <= data_in(5666);
     data_out(2435) <= data_in(5668);
     data_out(2436) <= data_in(5669);
     data_out(2437) <= data_in(5670);
     data_out(2438) <= data_in(5671);
     data_out(2439) <= data_in(5674);
     data_out(2440) <= data_in(5676);
     data_out(2441) <= data_in(5677);
     data_out(2442) <= data_in(5682);
     data_out(2443) <= data_in(5687);
     data_out(2444) <= data_in(5688);
     data_out(2445) <= data_in(5690);
     data_out(2446) <= data_in(5692);
     data_out(2447) <= data_in(5695);
     data_out(2448) <= data_in(5697);
     data_out(2449) <= data_in(5698);
     data_out(2450) <= data_in(5701);
     data_out(2451) <= data_in(5703);
     data_out(2452) <= data_in(5704);
     data_out(2453) <= data_in(5705);
     data_out(2454) <= data_in(5707);
     data_out(2455) <= data_in(5708);
     data_out(2456) <= data_in(5710);
     data_out(2457) <= data_in(5715);
     data_out(2458) <= data_in(5716);
     data_out(2459) <= data_in(5717);
     data_out(2460) <= data_in(5718);
     data_out(2461) <= data_in(5722);
     data_out(2462) <= data_in(5725);
     data_out(2463) <= data_in(5727);
     data_out(2464) <= data_in(5728);
     data_out(2465) <= data_in(5729);
     data_out(2466) <= data_in(5731);
     data_out(2467) <= data_in(5734);
     data_out(2468) <= data_in(5735);
     data_out(2469) <= data_in(5738);
     data_out(2470) <= data_in(5739);
     data_out(2471) <= data_in(5746);
     data_out(2472) <= data_in(5748);
     data_out(2473) <= data_in(5751);
     data_out(2474) <= data_in(5756);
     data_out(2475) <= data_in(5758);
     data_out(2476) <= data_in(5760);
     data_out(2477) <= data_in(5762);
     data_out(2478) <= data_in(5763);
     data_out(2479) <= data_in(5766);
     data_out(2480) <= data_in(5770);
     data_out(2481) <= data_in(5771);
     data_out(2482) <= data_in(5773);
     data_out(2483) <= data_in(5775);
     data_out(2484) <= data_in(5780);
     data_out(2485) <= data_in(5781);
     data_out(2486) <= data_in(5784);
     data_out(2487) <= data_in(5787);
     data_out(2488) <= data_in(5788);
     data_out(2489) <= data_in(5789);
     data_out(2490) <= data_in(5792);
     data_out(2491) <= data_in(5796);
     data_out(2492) <= data_in(5798);
     data_out(2493) <= data_in(5799);
     data_out(2494) <= data_in(5808);
     data_out(2495) <= data_in(5811);
     data_out(2496) <= data_in(5812);
     data_out(2497) <= data_in(5813);
     data_out(2498) <= data_in(5818);
     data_out(2499) <= data_in(5820);
     data_out(2500) <= data_in(5821);
     data_out(2501) <= data_in(5822);
     data_out(2502) <= data_in(5826);
     data_out(2503) <= data_in(5827);
     data_out(2504) <= data_in(5828);
     data_out(2505) <= data_in(5830);
     data_out(2506) <= data_in(5833);
     data_out(2507) <= data_in(5834);
     data_out(2508) <= data_in(5836);
     data_out(2509) <= data_in(5837);
     data_out(2510) <= data_in(5839);
     data_out(2511) <= data_in(5845);
     data_out(2512) <= data_in(5847);
     data_out(2513) <= data_in(5851);
     data_out(2514) <= data_in(5853);
     data_out(2515) <= data_in(5854);
     data_out(2516) <= data_in(5855);
     data_out(2517) <= data_in(5857);
     data_out(2518) <= data_in(5859);
     data_out(2519) <= data_in(5868);
     data_out(2520) <= data_in(5869);
     data_out(2521) <= data_in(5873);
     data_out(2522) <= data_in(5875);
     data_out(2523) <= data_in(5877);
     data_out(2524) <= data_in(5878);
     data_out(2525) <= data_in(5882);
     data_out(2526) <= data_in(5884);
     data_out(2527) <= data_in(5886);
     data_out(2528) <= data_in(5888);
     data_out(2529) <= data_in(5889);
     data_out(2530) <= data_in(5891);
     data_out(2531) <= data_in(5892);
     data_out(2532) <= data_in(5893);
     data_out(2533) <= data_in(5895);
     data_out(2534) <= data_in(5896);
     data_out(2535) <= data_in(5897);
     data_out(2536) <= data_in(5900);
     data_out(2537) <= data_in(5904);
     data_out(2538) <= data_in(5911);
     data_out(2539) <= data_in(5913);
     data_out(2540) <= data_in(5915);
     data_out(2541) <= data_in(5916);
     data_out(2542) <= data_in(5917);
     data_out(2543) <= data_in(5918);
     data_out(2544) <= data_in(5920);
     data_out(2545) <= data_in(5926);
     data_out(2546) <= data_in(5927);
     data_out(2547) <= data_in(5936);
     data_out(2548) <= data_in(5939);
     data_out(2549) <= data_in(5940);
     data_out(2550) <= data_in(5941);
     data_out(2551) <= data_in(5944);
     data_out(2552) <= data_in(5946);
     data_out(2553) <= data_in(5947);
     data_out(2554) <= data_in(5948);
     data_out(2555) <= data_in(5949);
     data_out(2556) <= data_in(5951);
     data_out(2557) <= data_in(5952);
     data_out(2558) <= data_in(5955);
     data_out(2559) <= data_in(5957);
     data_out(2560) <= data_in(5962);
     data_out(2561) <= data_in(5968);
     data_out(2562) <= data_in(5969);
     data_out(2563) <= data_in(5970);
     data_out(2564) <= data_in(5972);
     data_out(2565) <= data_in(5977);
     data_out(2566) <= data_in(5978);
     data_out(2567) <= data_in(5980);
     data_out(2568) <= data_in(5982);
     data_out(2569) <= data_in(5990);
     data_out(2570) <= data_in(5991);
     data_out(2571) <= data_in(5993);
     data_out(2572) <= data_in(5994);
     data_out(2573) <= data_in(5995);
     data_out(2574) <= data_in(6000);
     data_out(2575) <= data_in(6001);
     data_out(2576) <= data_in(6004);
     data_out(2577) <= data_in(6007);
     data_out(2578) <= data_in(6008);
     data_out(2579) <= data_in(6009);
     data_out(2580) <= data_in(6010);
     data_out(2581) <= data_in(6012);
     data_out(2582) <= data_in(6023);
     data_out(2583) <= data_in(6024);
     data_out(2584) <= data_in(6027);
     data_out(2585) <= data_in(6028);
     data_out(2586) <= data_in(6030);
     data_out(2587) <= data_in(6032);
     data_out(2588) <= data_in(6033);
     data_out(2589) <= data_in(6036);
     data_out(2590) <= data_in(6038);
     data_out(2591) <= data_in(6040);
     data_out(2592) <= data_in(6041);
     data_out(2593) <= data_in(6050);
     data_out(2594) <= data_in(6051);
     data_out(2595) <= data_in(6056);
     data_out(2596) <= data_in(6058);
     data_out(2597) <= data_in(6062);
     data_out(2598) <= data_in(6064);
     data_out(2599) <= data_in(6066);
     data_out(2600) <= data_in(6067);
     data_out(2601) <= data_in(6068);
     data_out(2602) <= data_in(6070);
     data_out(2603) <= data_in(6074);
     data_out(2604) <= data_in(6075);
     data_out(2605) <= data_in(6078);
     data_out(2606) <= data_in(6079);
     data_out(2607) <= data_in(6081);
     data_out(2608) <= data_in(6085);
     data_out(2609) <= data_in(6088);
     data_out(2610) <= data_in(6090);
     data_out(2611) <= data_in(6097);
     data_out(2612) <= data_in(6106);
     data_out(2613) <= data_in(6110);
     data_out(2614) <= data_in(6111);
     data_out(2615) <= data_in(6115);
     data_out(2616) <= data_in(6116);
     data_out(2617) <= data_in(6119);
     data_out(2618) <= data_in(6120);
     data_out(2619) <= data_in(6122);
     data_out(2620) <= data_in(6123);
     data_out(2621) <= data_in(6126);
     data_out(2622) <= data_in(6128);
     data_out(2623) <= data_in(6129);
     data_out(2624) <= data_in(6131);
     data_out(2625) <= data_in(6132);
     data_out(2626) <= data_in(6136);
     data_out(2627) <= data_in(6137);
     data_out(2628) <= data_in(6138);
     data_out(2629) <= data_in(6139);
     data_out(2630) <= data_in(6140);
     data_out(2631) <= data_in(6144);
     data_out(2632) <= data_in(6145);
     data_out(2633) <= data_in(6148);
     data_out(2634) <= data_in(6151);
     data_out(2635) <= data_in(6152);
     data_out(2636) <= data_in(6157);
     data_out(2637) <= data_in(6160);
     data_out(2638) <= data_in(6168);
     data_out(2639) <= data_in(6170);
     data_out(2640) <= data_in(6172);
     data_out(2641) <= data_in(6173);
     data_out(2642) <= data_in(6175);
     data_out(2643) <= data_in(6176);
     data_out(2644) <= data_in(6178);
     data_out(2645) <= data_in(6181);
     data_out(2646) <= data_in(6182);
     data_out(2647) <= data_in(6184);
     data_out(2648) <= data_in(6192);
     data_out(2649) <= data_in(6194);
     data_out(2650) <= data_in(6197);
     data_out(2651) <= data_in(6198);
     data_out(2652) <= data_in(6204);
     data_out(2653) <= data_in(6206);
     data_out(2654) <= data_in(6207);
     data_out(2655) <= data_in(6208);
     data_out(2656) <= data_in(6210);
     data_out(2657) <= data_in(6214);
     data_out(2658) <= data_in(6215);
     data_out(2659) <= data_in(6216);
     data_out(2660) <= data_in(6217);
     data_out(2661) <= data_in(6218);
     data_out(2662) <= data_in(6221);
     data_out(2663) <= data_in(6223);
     data_out(2664) <= data_in(6225);
     data_out(2665) <= data_in(6226);
     data_out(2666) <= data_in(6234);
     data_out(2667) <= data_in(6237);
     data_out(2668) <= data_in(6238);
     data_out(2669) <= data_in(6239);
     data_out(2670) <= data_in(6242);
     data_out(2671) <= data_in(6249);
     data_out(2672) <= data_in(6250);
     data_out(2673) <= data_in(6251);
     data_out(2674) <= data_in(6252);
     data_out(2675) <= data_in(6253);
     data_out(2676) <= data_in(6255);
     data_out(2677) <= data_in(6256);
     data_out(2678) <= data_in(6261);
     data_out(2679) <= data_in(6263);
     data_out(2680) <= data_in(6265);
     data_out(2681) <= data_in(6269);
     data_out(2682) <= data_in(6273);
     data_out(2683) <= data_in(6274);
     data_out(2684) <= data_in(6276);
     data_out(2685) <= data_in(6280);
     data_out(2686) <= data_in(6286);
     data_out(2687) <= data_in(6289);
     data_out(2688) <= data_in(6291);
     data_out(2689) <= data_in(6293);
     data_out(2690) <= data_in(6294);
     data_out(2691) <= data_in(6296);
     data_out(2692) <= data_in(6301);
     data_out(2693) <= data_in(6302);
     data_out(2694) <= data_in(6306);
     data_out(2695) <= data_in(6308);
     data_out(2696) <= data_in(6310);
     data_out(2697) <= data_in(6316);
     data_out(2698) <= data_in(6321);
     data_out(2699) <= data_in(6322);
     data_out(2700) <= data_in(6326);
     data_out(2701) <= data_in(6327);
     data_out(2702) <= data_in(6330);
     data_out(2703) <= data_in(6335);
     data_out(2704) <= data_in(6338);
     data_out(2705) <= data_in(6342);
     data_out(2706) <= data_in(6343);
     data_out(2707) <= data_in(6344);
     data_out(2708) <= data_in(6346);
     data_out(2709) <= data_in(6349);
     data_out(2710) <= data_in(6351);
     data_out(2711) <= data_in(6355);
     data_out(2712) <= data_in(6356);
     data_out(2713) <= data_in(6357);
     data_out(2714) <= data_in(6358);
     data_out(2715) <= data_in(6361);
     data_out(2716) <= data_in(6363);
     data_out(2717) <= data_in(6365);
     data_out(2718) <= data_in(6367);
     data_out(2719) <= data_in(6368);
     data_out(2720) <= data_in(6370);
     data_out(2721) <= data_in(6374);
     data_out(2722) <= data_in(6378);
     data_out(2723) <= data_in(6381);
     data_out(2724) <= data_in(6384);
     data_out(2725) <= data_in(6385);
     data_out(2726) <= data_in(6388);
     data_out(2727) <= data_in(6390);
     data_out(2728) <= data_in(6391);
     data_out(2729) <= data_in(6392);
     data_out(2730) <= data_in(6393);
     data_out(2731) <= data_in(6394);
     data_out(2732) <= data_in(6398);
     data_out(2733) <= data_in(6399);
     data_out(2734) <= data_in(6401);
     data_out(2735) <= data_in(6402);
     data_out(2736) <= data_in(6404);
     data_out(2737) <= data_in(6406);
     data_out(2738) <= data_in(6410);
     data_out(2739) <= data_in(6416);
     data_out(2740) <= data_in(6418);
     data_out(2741) <= data_in(6422);
     data_out(2742) <= data_in(6424);
     data_out(2743) <= data_in(6426);
     data_out(2744) <= data_in(6434);
     data_out(2745) <= data_in(6435);
     data_out(2746) <= data_in(6439);
     data_out(2747) <= data_in(6443);
     data_out(2748) <= data_in(6444);
     data_out(2749) <= data_in(6446);
     data_out(2750) <= data_in(6449);
     data_out(2751) <= data_in(6451);
     data_out(2752) <= data_in(6456);
     data_out(2753) <= data_in(6461);
     data_out(2754) <= data_in(6464);
     data_out(2755) <= data_in(6466);
     data_out(2756) <= data_in(6468);
     data_out(2757) <= data_in(6470);
     data_out(2758) <= data_in(6473);
     data_out(2759) <= data_in(6481);
     data_out(2760) <= data_in(6482);
     data_out(2761) <= data_in(6483);
     data_out(2762) <= data_in(6486);
     data_out(2763) <= data_in(6488);
     data_out(2764) <= data_in(6489);
     data_out(2765) <= data_in(6490);
     data_out(2766) <= data_in(6491);
     data_out(2767) <= data_in(6492);
     data_out(2768) <= data_in(6493);
     data_out(2769) <= data_in(6494);
     data_out(2770) <= data_in(6495);
     data_out(2771) <= data_in(6496);
     data_out(2772) <= data_in(6497);
     data_out(2773) <= data_in(6504);
     data_out(2774) <= data_in(6509);
     data_out(2775) <= data_in(6511);
     data_out(2776) <= data_in(6513);
     data_out(2777) <= data_in(6514);
     data_out(2778) <= data_in(6519);
     data_out(2779) <= data_in(6521);
     data_out(2780) <= data_in(6522);
     data_out(2781) <= data_in(6528);
     data_out(2782) <= data_in(6531);
     data_out(2783) <= data_in(6533);
     data_out(2784) <= data_in(6536);
     data_out(2785) <= data_in(6537);
     data_out(2786) <= data_in(6538);
     data_out(2787) <= data_in(6539);
     data_out(2788) <= data_in(6540);
     data_out(2789) <= data_in(6541);
     data_out(2790) <= data_in(6542);
     data_out(2791) <= data_in(6545);
     data_out(2792) <= data_in(6547);
     data_out(2793) <= data_in(6550);
     data_out(2794) <= data_in(6552);
     data_out(2795) <= data_in(6554);
     data_out(2796) <= data_in(6556);
     data_out(2797) <= data_in(6557);
     data_out(2798) <= data_in(6559);
     data_out(2799) <= data_in(6560);
     data_out(2800) <= data_in(6562);
     data_out(2801) <= data_in(6568);
     data_out(2802) <= data_in(6569);
     data_out(2803) <= data_in(6574);
     data_out(2804) <= data_in(6575);
     data_out(2805) <= data_in(6576);
     data_out(2806) <= data_in(6579);
     data_out(2807) <= data_in(6580);
     data_out(2808) <= data_in(6581);
     data_out(2809) <= data_in(6582);
     data_out(2810) <= data_in(6586);
     data_out(2811) <= data_in(6589);
     data_out(2812) <= data_in(6590);
     data_out(2813) <= data_in(6591);
     data_out(2814) <= data_in(6594);
     data_out(2815) <= data_in(6601);
     data_out(2816) <= data_in(6603);
     data_out(2817) <= data_in(6604);
     data_out(2818) <= data_in(6606);
     data_out(2819) <= data_in(6607);
     data_out(2820) <= data_in(6608);
     data_out(2821) <= data_in(6609);
     data_out(2822) <= data_in(6610);
     data_out(2823) <= data_in(6613);
     data_out(2824) <= data_in(6616);
     data_out(2825) <= data_in(6619);
     data_out(2826) <= data_in(6620);
     data_out(2827) <= data_in(6624);
     data_out(2828) <= data_in(6625);
     data_out(2829) <= data_in(6628);
     data_out(2830) <= data_in(6629);
     data_out(2831) <= data_in(6634);
     data_out(2832) <= data_in(6635);
     data_out(2833) <= data_in(6638);
     data_out(2834) <= data_in(6641);
     data_out(2835) <= data_in(6642);
     data_out(2836) <= data_in(6643);
     data_out(2837) <= data_in(6648);
     data_out(2838) <= data_in(6649);
     data_out(2839) <= data_in(6650);
     data_out(2840) <= data_in(6651);
     data_out(2841) <= data_in(6654);
     data_out(2842) <= data_in(6657);
     data_out(2843) <= data_in(6658);
     data_out(2844) <= data_in(6660);
     data_out(2845) <= data_in(6661);
     data_out(2846) <= data_in(6665);
     data_out(2847) <= data_in(6668);
     data_out(2848) <= data_in(6670);
     data_out(2849) <= data_in(6671);
     data_out(2850) <= data_in(6675);
     data_out(2851) <= data_in(6677);
     data_out(2852) <= data_in(6679);
     data_out(2853) <= data_in(6680);
     data_out(2854) <= data_in(6681);
     data_out(2855) <= data_in(6684);
     data_out(2856) <= data_in(6686);
     data_out(2857) <= data_in(6693);
     data_out(2858) <= data_in(6694);
     data_out(2859) <= data_in(6695);
     data_out(2860) <= data_in(6696);
     data_out(2861) <= data_in(6699);
     data_out(2862) <= data_in(6702);
     data_out(2863) <= data_in(6703);
     data_out(2864) <= data_in(6704);
     data_out(2865) <= data_in(6705);
     data_out(2866) <= data_in(6706);
     data_out(2867) <= data_in(6707);
     data_out(2868) <= data_in(6708);
     data_out(2869) <= data_in(6709);
     data_out(2870) <= data_in(6710);
     data_out(2871) <= data_in(6711);
     data_out(2872) <= data_in(6720);
     data_out(2873) <= data_in(6724);
     data_out(2874) <= data_in(6726);
     data_out(2875) <= data_in(6727);
     data_out(2876) <= data_in(6728);
     data_out(2877) <= data_in(6730);
     data_out(2878) <= data_in(6738);
     data_out(2879) <= data_in(6740);
     data_out(2880) <= data_in(6742);
     data_out(2881) <= data_in(6744);
     data_out(2882) <= data_in(6745);
     data_out(2883) <= data_in(6746);
     data_out(2884) <= data_in(6748);
     data_out(2885) <= data_in(6753);
     data_out(2886) <= data_in(6755);
     data_out(2887) <= data_in(6757);
     data_out(2888) <= data_in(6760);
     data_out(2889) <= data_in(6761);
     data_out(2890) <= data_in(6762);
     data_out(2891) <= data_in(6763);
     data_out(2892) <= data_in(6768);
     data_out(2893) <= data_in(6773);
     data_out(2894) <= data_in(6774);
     data_out(2895) <= data_in(6780);
     data_out(2896) <= data_in(6782);
     data_out(2897) <= data_in(6785);
     data_out(2898) <= data_in(6786);
     data_out(2899) <= data_in(6787);
     data_out(2900) <= data_in(6788);
     data_out(2901) <= data_in(6791);
     data_out(2902) <= data_in(6793);
     data_out(2903) <= data_in(6794);
     data_out(2904) <= data_in(6795);
     data_out(2905) <= data_in(6797);
     data_out(2906) <= data_in(6804);
     data_out(2907) <= data_in(6805);
     data_out(2908) <= data_in(6806);
     data_out(2909) <= data_in(6807);
     data_out(2910) <= data_in(6809);
     data_out(2911) <= data_in(6812);
     data_out(2912) <= data_in(6817);
     data_out(2913) <= data_in(6818);
     data_out(2914) <= data_in(6820);
     data_out(2915) <= data_in(6821);
     data_out(2916) <= data_in(6823);
     data_out(2917) <= data_in(6825);
     data_out(2918) <= data_in(6826);
     data_out(2919) <= data_in(6827);
     data_out(2920) <= data_in(6834);
     data_out(2921) <= data_in(6838);
     data_out(2922) <= data_in(6840);
     data_out(2923) <= data_in(6842);
     data_out(2924) <= data_in(6844);
     data_out(2925) <= data_in(6845);
     data_out(2926) <= data_in(6846);
     data_out(2927) <= data_in(6848);
     data_out(2928) <= data_in(6849);
     data_out(2929) <= data_in(6853);
     data_out(2930) <= data_in(6855);
     data_out(2931) <= data_in(6857);
     data_out(2932) <= data_in(6859);
     data_out(2933) <= data_in(6862);
     data_out(2934) <= data_in(6863);
     data_out(2935) <= data_in(6864);
     data_out(2936) <= data_in(6867);
     data_out(2937) <= data_in(6868);
     data_out(2938) <= data_in(6869);
     data_out(2939) <= data_in(6870);
     data_out(2940) <= data_in(6871);
     data_out(2941) <= data_in(6879);
     data_out(2942) <= data_in(6880);
     data_out(2943) <= data_in(6881);
     data_out(2944) <= data_in(6882);
     data_out(2945) <= data_in(6883);
     data_out(2946) <= data_in(6885);
     data_out(2947) <= data_in(6888);
     data_out(2948) <= data_in(6890);
     data_out(2949) <= data_in(6892);
     data_out(2950) <= data_in(6894);
     data_out(2951) <= data_in(6895);
     data_out(2952) <= data_in(6896);
     data_out(2953) <= data_in(6897);
     data_out(2954) <= data_in(6901);
     data_out(2955) <= data_in(6902);
     data_out(2956) <= data_in(6905);
     data_out(2957) <= data_in(6907);
     data_out(2958) <= data_in(6909);
     data_out(2959) <= data_in(6913);
     data_out(2960) <= data_in(6917);
     data_out(2961) <= data_in(6920);
     data_out(2962) <= data_in(6922);
     data_out(2963) <= data_in(6924);
     data_out(2964) <= data_in(6925);
     data_out(2965) <= data_in(6926);
     data_out(2966) <= data_in(6927);
     data_out(2967) <= data_in(6928);
     data_out(2968) <= data_in(6929);
     data_out(2969) <= data_in(6933);
     data_out(2970) <= data_in(6937);
     data_out(2971) <= data_in(6939);
     data_out(2972) <= data_in(6941);
     data_out(2973) <= data_in(6942);
     data_out(2974) <= data_in(6943);
     data_out(2975) <= data_in(6947);
     data_out(2976) <= data_in(6949);
     data_out(2977) <= data_in(6950);
     data_out(2978) <= data_in(6952);
     data_out(2979) <= data_in(6957);
     data_out(2980) <= data_in(6958);
     data_out(2981) <= data_in(6959);
     data_out(2982) <= data_in(6961);
     data_out(2983) <= data_in(6962);
     data_out(2984) <= data_in(6967);
     data_out(2985) <= data_in(6969);
     data_out(2986) <= data_in(6971);
     data_out(2987) <= data_in(6972);
     data_out(2988) <= data_in(6974);
     data_out(2989) <= data_in(6976);
     data_out(2990) <= data_in(6978);
     data_out(2991) <= data_in(6979);
     data_out(2992) <= data_in(6980);
     data_out(2993) <= data_in(6981);
     data_out(2994) <= data_in(6982);
     data_out(2995) <= data_in(6984);
     data_out(2996) <= data_in(6986);
     data_out(2997) <= data_in(6989);
     data_out(2998) <= data_in(6990);
     data_out(2999) <= data_in(6997);
     data_out(3000) <= data_in(7002);
     data_out(3001) <= data_in(7003);
     data_out(3002) <= data_in(7006);
     data_out(3003) <= data_in(7010);
     data_out(3004) <= data_in(7012);
     data_out(3005) <= data_in(7015);
     data_out(3006) <= data_in(7016);
     data_out(3007) <= data_in(7017);
     data_out(3008) <= data_in(7019);
     data_out(3009) <= data_in(7022);
     data_out(3010) <= data_in(7023);
     data_out(3011) <= data_in(7025);
     data_out(3012) <= data_in(7026);
     data_out(3013) <= data_in(7030);
     data_out(3014) <= data_in(7035);
     data_out(3015) <= data_in(7036);
     data_out(3016) <= data_in(7038);
     data_out(3017) <= data_in(7039);
     data_out(3018) <= data_in(7041);
     data_out(3019) <= data_in(7042);
     data_out(3020) <= data_in(7043);
     data_out(3021) <= data_in(7044);
     data_out(3022) <= data_in(7046);
     data_out(3023) <= data_in(7047);
     data_out(3024) <= data_in(7048);
     data_out(3025) <= data_in(7049);
     data_out(3026) <= data_in(7058);
     data_out(3027) <= data_in(7060);
     data_out(3028) <= data_in(7064);
     data_out(3029) <= data_in(7065);
     data_out(3030) <= data_in(7068);
     data_out(3031) <= data_in(7070);
     data_out(3032) <= data_in(7080);
     data_out(3033) <= data_in(7081);
     data_out(3034) <= data_in(7082);
     data_out(3035) <= data_in(7083);
     data_out(3036) <= data_in(7089);
     data_out(3037) <= data_in(7091);
     data_out(3038) <= data_in(7097);
     data_out(3039) <= data_in(7099);
     data_out(3040) <= data_in(7101);
     data_out(3041) <= data_in(7104);
     data_out(3042) <= data_in(7106);
     data_out(3043) <= data_in(7108);
     data_out(3044) <= data_in(7110);
     data_out(3045) <= data_in(7111);
     data_out(3046) <= data_in(7113);
     data_out(3047) <= data_in(7114);
     data_out(3048) <= data_in(7116);
     data_out(3049) <= data_in(7117);
     data_out(3050) <= data_in(7118);
     data_out(3051) <= data_in(7122);
     data_out(3052) <= data_in(7124);
     data_out(3053) <= data_in(7127);
     data_out(3054) <= data_in(7128);
     data_out(3055) <= data_in(7129);
     data_out(3056) <= data_in(7133);
     data_out(3057) <= data_in(7134);
     data_out(3058) <= data_in(7137);
     data_out(3059) <= data_in(7138);
     data_out(3060) <= data_in(7139);
     data_out(3061) <= data_in(7140);
     data_out(3062) <= data_in(7142);
     data_out(3063) <= data_in(7143);
     data_out(3064) <= data_in(7144);
     data_out(3065) <= data_in(7147);
     data_out(3066) <= data_in(7150);
     data_out(3067) <= data_in(7151);
     data_out(3068) <= data_in(7154);
     data_out(3069) <= data_in(7157);
     data_out(3070) <= data_in(7159);
     data_out(3071) <= data_in(7162);
     data_out(3072) <= data_in(7164);
     data_out(3073) <= data_in(7165);
     data_out(3074) <= data_in(7171);
     data_out(3075) <= data_in(7173);
     data_out(3076) <= data_in(7178);
     data_out(3077) <= data_in(7181);
     data_out(3078) <= data_in(7185);
     data_out(3079) <= data_in(7189);
     data_out(3080) <= data_in(7190);
     data_out(3081) <= data_in(7193);
     data_out(3082) <= data_in(7195);
     data_out(3083) <= data_in(7197);
     data_out(3084) <= data_in(7202);
     data_out(3085) <= data_in(7204);
     data_out(3086) <= data_in(7206);
     data_out(3087) <= data_in(7210);
     data_out(3088) <= data_in(7212);
     data_out(3089) <= data_in(7213);
     data_out(3090) <= data_in(7214);
     data_out(3091) <= data_in(7215);
     data_out(3092) <= data_in(7219);
     data_out(3093) <= data_in(7224);
     data_out(3094) <= data_in(7226);
     data_out(3095) <= data_in(7228);
     data_out(3096) <= data_in(7230);
     data_out(3097) <= data_in(7231);
     data_out(3098) <= data_in(7233);
     data_out(3099) <= data_in(7236);
     data_out(3100) <= data_in(7240);
     data_out(3101) <= data_in(7246);
     data_out(3102) <= data_in(7248);
     data_out(3103) <= data_in(7249);
     data_out(3104) <= data_in(7256);
     data_out(3105) <= data_in(7257);
     data_out(3106) <= data_in(7262);
     data_out(3107) <= data_in(7270);
     data_out(3108) <= data_in(7273);
     data_out(3109) <= data_in(7275);
     data_out(3110) <= data_in(7277);
     data_out(3111) <= data_in(7285);
     data_out(3112) <= data_in(7291);
     data_out(3113) <= data_in(7292);
     data_out(3114) <= data_in(7296);
     data_out(3115) <= data_in(7297);
     data_out(3116) <= data_in(7298);
     data_out(3117) <= data_in(7299);
     data_out(3118) <= data_in(7300);
     data_out(3119) <= data_in(7304);
     data_out(3120) <= data_in(7307);
     data_out(3121) <= data_in(7309);
     data_out(3122) <= data_in(7311);
     data_out(3123) <= data_in(7315);
     data_out(3124) <= data_in(7321);
     data_out(3125) <= data_in(7322);
     data_out(3126) <= data_in(7327);
     data_out(3127) <= data_in(7330);
     data_out(3128) <= data_in(7333);
     data_out(3129) <= data_in(7334);
     data_out(3130) <= data_in(7335);
     data_out(3131) <= data_in(7338);
     data_out(3132) <= data_in(7342);
     data_out(3133) <= data_in(7343);
     data_out(3134) <= data_in(7345);
     data_out(3135) <= data_in(7346);
     data_out(3136) <= data_in(7347);
     data_out(3137) <= data_in(7349);
     data_out(3138) <= data_in(7350);
     data_out(3139) <= data_in(7351);
     data_out(3140) <= data_in(7352);
     data_out(3141) <= data_in(7354);
     data_out(3142) <= data_in(7356);
     data_out(3143) <= data_in(7357);
     data_out(3144) <= data_in(7360);
     data_out(3145) <= data_in(7361);
     data_out(3146) <= data_in(7363);
     data_out(3147) <= data_in(7368);
     data_out(3148) <= data_in(7370);
     data_out(3149) <= data_in(7371);
     data_out(3150) <= data_in(7372);
     data_out(3151) <= data_in(7376);
     data_out(3152) <= data_in(7378);
     data_out(3153) <= data_in(7385);
     data_out(3154) <= data_in(7387);
     data_out(3155) <= data_in(7390);
     data_out(3156) <= data_in(7391);
     data_out(3157) <= data_in(7393);
     data_out(3158) <= data_in(7394);
     data_out(3159) <= data_in(7397);
     data_out(3160) <= data_in(7398);
     data_out(3161) <= data_in(7399);
     data_out(3162) <= data_in(7401);
     data_out(3163) <= data_in(7404);
     data_out(3164) <= data_in(7408);
     data_out(3165) <= data_in(7411);
     data_out(3166) <= data_in(7414);
     data_out(3167) <= data_in(7417);
     data_out(3168) <= data_in(7425);
     data_out(3169) <= data_in(7426);
     data_out(3170) <= data_in(7432);
     data_out(3171) <= data_in(7435);
     data_out(3172) <= data_in(7436);
     data_out(3173) <= data_in(7441);
     data_out(3174) <= data_in(7442);
     data_out(3175) <= data_in(7443);
     data_out(3176) <= data_in(7446);
     data_out(3177) <= data_in(7450);
     data_out(3178) <= data_in(7451);
     data_out(3179) <= data_in(7452);
     data_out(3180) <= data_in(7454);
     data_out(3181) <= data_in(7455);
     data_out(3182) <= data_in(7465);
     data_out(3183) <= data_in(7466);
     data_out(3184) <= data_in(7467);
     data_out(3185) <= data_in(7468);
     data_out(3186) <= data_in(7469);
     data_out(3187) <= data_in(7471);
     data_out(3188) <= data_in(7474);
     data_out(3189) <= data_in(7475);
     data_out(3190) <= data_in(7479);
     data_out(3191) <= data_in(7480);
     data_out(3192) <= data_in(7481);
     data_out(3193) <= data_in(7483);
     data_out(3194) <= data_in(7484);
     data_out(3195) <= data_in(7487);
     data_out(3196) <= data_in(7489);
     data_out(3197) <= data_in(7495);
     data_out(3198) <= data_in(7496);
     data_out(3199) <= data_in(7499);
     data_out(3200) <= data_in(7500);
     data_out(3201) <= data_in(7501);
     data_out(3202) <= data_in(7502);
     data_out(3203) <= data_in(7504);
     data_out(3204) <= data_in(7517);
     data_out(3205) <= data_in(7519);
     data_out(3206) <= data_in(7520);
     data_out(3207) <= data_in(7521);
     data_out(3208) <= data_in(7525);
     data_out(3209) <= data_in(7528);
     data_out(3210) <= data_in(7530);
     data_out(3211) <= data_in(7531);
     data_out(3212) <= data_in(7535);
     data_out(3213) <= data_in(7537);
     data_out(3214) <= data_in(7539);
     data_out(3215) <= data_in(7541);
     data_out(3216) <= data_in(7542);
     data_out(3217) <= data_in(7543);
     data_out(3218) <= data_in(7547);
     data_out(3219) <= data_in(7548);
     data_out(3220) <= data_in(7549);
     data_out(3221) <= data_in(7551);
     data_out(3222) <= data_in(7552);
     data_out(3223) <= data_in(7554);
     data_out(3224) <= data_in(7571);
     data_out(3225) <= data_in(7573);
     data_out(3226) <= data_in(7575);
     data_out(3227) <= data_in(7576);
     data_out(3228) <= data_in(7577);
     data_out(3229) <= data_in(7578);
     data_out(3230) <= data_in(7579);
     data_out(3231) <= data_in(7584);
     data_out(3232) <= data_in(7586);
     data_out(3233) <= data_in(7587);
     data_out(3234) <= data_in(7589);
     data_out(3235) <= data_in(7592);
     data_out(3236) <= data_in(7593);
     data_out(3237) <= data_in(7594);
     data_out(3238) <= data_in(7595);
     data_out(3239) <= data_in(7597);
     data_out(3240) <= data_in(7598);
     data_out(3241) <= data_in(7599);
     data_out(3242) <= data_in(7602);
     data_out(3243) <= data_in(7606);
     data_out(3244) <= data_in(7607);
     data_out(3245) <= data_in(7609);
     data_out(3246) <= data_in(7612);
     data_out(3247) <= data_in(7613);
     data_out(3248) <= data_in(7614);
     data_out(3249) <= data_in(7615);
     data_out(3250) <= data_in(7621);
     data_out(3251) <= data_in(7622);
     data_out(3252) <= data_in(7623);
     data_out(3253) <= data_in(7624);
     data_out(3254) <= data_in(7625);
     data_out(3255) <= data_in(7626);
     data_out(3256) <= data_in(7643);
     data_out(3257) <= data_in(7644);
     data_out(3258) <= data_in(7646);
     data_out(3259) <= data_in(7647);
     data_out(3260) <= data_in(7648);
     data_out(3261) <= data_in(7654);
     data_out(3262) <= data_in(7661);
     data_out(3263) <= data_in(7666);
     data_out(3264) <= data_in(7672);
     data_out(3265) <= data_in(7677);
     data_out(3266) <= data_in(7678);
     data_out(3267) <= data_in(7679);
     data_out(3268) <= data_in(7680);
     data_out(3269) <= data_in(7681);
     data_out(3270) <= data_in(7686);
     data_out(3271) <= data_in(7688);
     data_out(3272) <= data_in(7690);
     data_out(3273) <= data_in(7693);
     data_out(3274) <= data_in(7694);
     data_out(3275) <= data_in(7695);
     data_out(3276) <= data_in(7698);
     data_out(3277) <= data_in(7699);
     data_out(3278) <= data_in(7701);
     data_out(3279) <= data_in(7704);
     data_out(3280) <= data_in(7705);
     data_out(3281) <= data_in(7706);
     data_out(3282) <= data_in(7707);
     data_out(3283) <= data_in(7714);
     data_out(3284) <= data_in(7717);
     data_out(3285) <= data_in(7721);
     data_out(3286) <= data_in(7724);
     data_out(3287) <= data_in(7726);
     data_out(3288) <= data_in(7727);
     data_out(3289) <= data_in(7728);
     data_out(3290) <= data_in(7730);
     data_out(3291) <= data_in(7737);
     data_out(3292) <= data_in(7739);
     data_out(3293) <= data_in(7740);
     data_out(3294) <= data_in(7743);
     data_out(3295) <= data_in(7744);
     data_out(3296) <= data_in(7746);
     data_out(3297) <= data_in(7749);
     data_out(3298) <= data_in(7759);
     data_out(3299) <= data_in(7760);
     data_out(3300) <= data_in(7762);
     data_out(3301) <= data_in(7764);
     data_out(3302) <= data_in(7769);
     data_out(3303) <= data_in(7771);
     data_out(3304) <= data_in(7774);
     data_out(3305) <= data_in(7775);
     data_out(3306) <= data_in(7777);
     data_out(3307) <= data_in(7778);
     data_out(3308) <= data_in(7779);
     data_out(3309) <= data_in(7781);
     data_out(3310) <= data_in(7782);
     data_out(3311) <= data_in(7784);
     data_out(3312) <= data_in(7792);
     data_out(3313) <= data_in(7793);
     data_out(3314) <= data_in(7798);
     data_out(3315) <= data_in(7800);
     data_out(3316) <= data_in(7803);
     data_out(3317) <= data_in(7804);
     data_out(3318) <= data_in(7808);
     data_out(3319) <= data_in(7809);
     data_out(3320) <= data_in(7810);
     data_out(3321) <= data_in(7814);
     data_out(3322) <= data_in(7815);
     data_out(3323) <= data_in(7819);
     data_out(3324) <= data_in(7823);
     data_out(3325) <= data_in(7824);
     data_out(3326) <= data_in(7825);
     data_out(3327) <= data_in(7826);
     data_out(3328) <= data_in(7827);
     data_out(3329) <= data_in(7833);
     data_out(3330) <= data_in(7835);
     data_out(3331) <= data_in(7836);
     data_out(3332) <= data_in(7838);
     data_out(3333) <= data_in(7849);
     data_out(3334) <= data_in(7850);
     data_out(3335) <= data_in(7851);
     data_out(3336) <= data_in(7852);
     data_out(3337) <= data_in(7854);
     data_out(3338) <= data_in(7855);
     data_out(3339) <= data_in(7859);
     data_out(3340) <= data_in(7860);
     data_out(3341) <= data_in(7862);
     data_out(3342) <= data_in(7864);
     data_out(3343) <= data_in(7869);
     data_out(3344) <= data_in(7870);
     data_out(3345) <= data_in(7872);
     data_out(3346) <= data_in(7874);
     data_out(3347) <= data_in(7875);
     data_out(3348) <= data_in(7879);
     data_out(3349) <= data_in(7880);
     data_out(3350) <= data_in(7881);
     data_out(3351) <= data_in(7882);
     data_out(3352) <= data_in(7883);
     data_out(3353) <= data_in(7884);
     data_out(3354) <= data_in(7886);
     data_out(3355) <= data_in(7889);
     data_out(3356) <= data_in(7893);
     data_out(3357) <= data_in(7894);
     data_out(3358) <= data_in(7897);
     data_out(3359) <= data_in(7898);
     data_out(3360) <= data_in(7900);
     data_out(3361) <= data_in(7907);
     data_out(3362) <= data_in(7908);
     data_out(3363) <= data_in(7909);
     data_out(3364) <= data_in(7910);
     data_out(3365) <= data_in(7917);
     data_out(3366) <= data_in(7918);
     data_out(3367) <= data_in(7922);
     data_out(3368) <= data_in(7924);
     data_out(3369) <= data_in(7926);
     data_out(3370) <= data_in(7927);
     data_out(3371) <= data_in(7937);
     data_out(3372) <= data_in(7939);
     data_out(3373) <= data_in(7945);
     data_out(3374) <= data_in(7948);
     data_out(3375) <= data_in(7952);
     data_out(3376) <= data_in(7953);
     data_out(3377) <= data_in(7960);
     data_out(3378) <= data_in(7961);
     data_out(3379) <= data_in(7963);
     data_out(3380) <= data_in(7964);
     data_out(3381) <= data_in(7969);
     data_out(3382) <= data_in(7970);
     data_out(3383) <= data_in(7971);
     data_out(3384) <= data_in(7977);
     data_out(3385) <= data_in(7980);
     data_out(3386) <= data_in(7983);
     data_out(3387) <= data_in(7984);
     data_out(3388) <= data_in(7986);
     data_out(3389) <= data_in(7989);
     data_out(3390) <= data_in(7993);
     data_out(3391) <= data_in(7994);
     data_out(3392) <= data_in(7995);
     data_out(3393) <= data_in(7996);
     data_out(3394) <= data_in(7997);
     data_out(3395) <= data_in(7998);
     data_out(3396) <= data_in(8002);
     data_out(3397) <= data_in(8005);
     data_out(3398) <= data_in(8008);
     data_out(3399) <= data_in(8010);
     data_out(3400) <= data_in(8012);
     data_out(3401) <= data_in(8014);
     data_out(3402) <= data_in(8019);
     data_out(3403) <= data_in(8022);
     data_out(3404) <= data_in(8031);
     data_out(3405) <= data_in(8033);
     data_out(3406) <= data_in(8035);
     data_out(3407) <= data_in(8036);
     data_out(3408) <= data_in(8038);
     data_out(3409) <= data_in(8039);
     data_out(3410) <= data_in(8042);
     data_out(3411) <= data_in(8043);
     data_out(3412) <= data_in(8044);
     data_out(3413) <= data_in(8045);
     data_out(3414) <= data_in(8046);
     data_out(3415) <= data_in(8051);
     data_out(3416) <= data_in(8052);
     data_out(3417) <= data_in(8054);
     data_out(3418) <= data_in(8055);
     data_out(3419) <= data_in(8056);
     data_out(3420) <= data_in(8059);
     data_out(3421) <= data_in(8060);
     data_out(3422) <= data_in(8062);
     data_out(3423) <= data_in(8064);
     data_out(3424) <= data_in(8066);
     data_out(3425) <= data_in(8067);
     data_out(3426) <= data_in(8068);
     data_out(3427) <= data_in(8070);
     data_out(3428) <= data_in(8072);
     data_out(3429) <= data_in(8078);
     data_out(3430) <= data_in(8079);
     data_out(3431) <= data_in(8081);
     data_out(3432) <= data_in(8082);
     data_out(3433) <= data_in(8084);
     data_out(3434) <= data_in(8085);
     data_out(3435) <= data_in(8087);
     data_out(3436) <= data_in(8093);
     data_out(3437) <= data_in(8095);
     data_out(3438) <= data_in(8096);
     data_out(3439) <= data_in(8097);
     data_out(3440) <= data_in(8102);
     data_out(3441) <= data_in(8115);
     data_out(3442) <= data_in(8124);
     data_out(3443) <= data_in(8127);
     data_out(3444) <= data_in(8130);
     data_out(3445) <= data_in(8132);
     data_out(3446) <= data_in(8139);
     data_out(3447) <= data_in(8140);
     data_out(3448) <= data_in(8141);
     data_out(3449) <= data_in(8142);
     data_out(3450) <= data_in(8143);
     data_out(3451) <= data_in(8144);
     data_out(3452) <= data_in(8148);
     data_out(3453) <= data_in(8149);
     data_out(3454) <= data_in(8150);
     data_out(3455) <= data_in(8158);
     data_out(3456) <= data_in(8159);
     data_out(3457) <= data_in(8164);
     data_out(3458) <= data_in(8166);
     data_out(3459) <= data_in(8167);
     data_out(3460) <= data_in(8169);
     data_out(3461) <= data_in(8172);
     data_out(3462) <= data_in(8178);
     data_out(3463) <= data_in(8179);
     data_out(3464) <= data_in(8180);
     data_out(3465) <= data_in(8182);
     data_out(3466) <= data_in(8188);
     data_out(3467) <= data_in(8194);
     data_out(3468) <= data_in(8196);
     data_out(3469) <= data_in(8199);
     data_out(3470) <= data_in(8201);
     data_out(3471) <= data_in(8208);
     data_out(3472) <= data_in(8209);
     data_out(3473) <= data_in(8211);
     data_out(3474) <= data_in(8214);
     data_out(3475) <= data_in(8215);
     data_out(3476) <= data_in(8216);
     data_out(3477) <= data_in(8220);
     data_out(3478) <= data_in(8224);
     data_out(3479) <= data_in(8225);
     data_out(3480) <= data_in(8227);
     data_out(3481) <= data_in(8229);
     data_out(3482) <= data_in(8232);
     data_out(3483) <= data_in(8236);
     data_out(3484) <= data_in(8239);
     data_out(3485) <= data_in(8240);
     data_out(3486) <= data_in(8246);
     data_out(3487) <= data_in(8247);
     data_out(3488) <= data_in(8248);
     data_out(3489) <= data_in(8249);
     data_out(3490) <= data_in(8250);
     data_out(3491) <= data_in(8254);
     data_out(3492) <= data_in(8260);
     data_out(3493) <= data_in(8261);
     data_out(3494) <= data_in(8264);
     data_out(3495) <= data_in(8265);
     data_out(3496) <= data_in(8269);
     data_out(3497) <= data_in(8272);
     data_out(3498) <= data_in(8274);
     data_out(3499) <= data_in(8275);
     data_out(3500) <= data_in(8276);
     data_out(3501) <= data_in(8280);
     data_out(3502) <= data_in(8284);
     data_out(3503) <= data_in(8289);
     data_out(3504) <= data_in(8290);
     data_out(3505) <= data_in(8291);
     data_out(3506) <= data_in(8292);
     data_out(3507) <= data_in(8293);
     data_out(3508) <= data_in(8295);
     data_out(3509) <= data_in(8296);
     data_out(3510) <= data_in(8305);
     data_out(3511) <= data_in(8310);
     data_out(3512) <= data_in(8317);
     data_out(3513) <= data_in(8319);
     data_out(3514) <= data_in(8320);
     data_out(3515) <= data_in(8323);
     data_out(3516) <= data_in(8326);
     data_out(3517) <= data_in(8329);
     data_out(3518) <= data_in(8330);
     data_out(3519) <= data_in(8331);
     data_out(3520) <= data_in(8333);
     data_out(3521) <= data_in(8334);
     data_out(3522) <= data_in(8336);
     data_out(3523) <= data_in(8340);
     data_out(3524) <= data_in(8341);
     data_out(3525) <= data_in(8342);
     data_out(3526) <= data_in(8343);
     data_out(3527) <= data_in(8345);
     data_out(3528) <= data_in(8347);
     data_out(3529) <= data_in(8353);
     data_out(3530) <= data_in(8355);
     data_out(3531) <= data_in(8356);
     data_out(3532) <= data_in(8361);
     data_out(3533) <= data_in(8364);
     data_out(3534) <= data_in(8367);
     data_out(3535) <= data_in(8368);
     data_out(3536) <= data_in(8375);
     data_out(3537) <= data_in(8376);
     data_out(3538) <= data_in(8377);
     data_out(3539) <= data_in(8381);
     data_out(3540) <= data_in(8382);
     data_out(3541) <= data_in(8388);
     data_out(3542) <= data_in(8392);
     data_out(3543) <= data_in(8394);
     data_out(3544) <= data_in(8400);
     data_out(3545) <= data_in(8402);
     data_out(3546) <= data_in(8403);
     data_out(3547) <= data_in(8406);
     data_out(3548) <= data_in(8407);
     data_out(3549) <= data_in(8408);
     data_out(3550) <= data_in(8409);
     data_out(3551) <= data_in(8412);
     data_out(3552) <= data_in(8413);
     data_out(3553) <= data_in(8417);
     data_out(3554) <= data_in(8420);
     data_out(3555) <= data_in(8421);
     data_out(3556) <= data_in(8422);
     data_out(3557) <= data_in(8425);
     data_out(3558) <= data_in(8428);
     data_out(3559) <= data_in(8430);
     data_out(3560) <= data_in(8431);
     data_out(3561) <= data_in(8433);
     data_out(3562) <= data_in(8437);
     data_out(3563) <= data_in(8439);
     data_out(3564) <= data_in(8440);
     data_out(3565) <= data_in(8441);
     data_out(3566) <= data_in(8443);
     data_out(3567) <= data_in(8444);
     data_out(3568) <= data_in(8446);
     data_out(3569) <= data_in(8450);
     data_out(3570) <= data_in(8452);
     data_out(3571) <= data_in(8453);
     data_out(3572) <= data_in(8457);
     data_out(3573) <= data_in(8458);
     data_out(3574) <= data_in(8459);
     data_out(3575) <= data_in(8460);
     data_out(3576) <= data_in(8462);
     data_out(3577) <= data_in(8468);
     data_out(3578) <= data_in(8469);
     data_out(3579) <= data_in(8470);
     data_out(3580) <= data_in(8471);
     data_out(3581) <= data_in(8473);
     data_out(3582) <= data_in(8476);
     data_out(3583) <= data_in(8477);
     data_out(3584) <= data_in(8479);
     data_out(3585) <= data_in(8482);
     data_out(3586) <= data_in(8484);
     data_out(3587) <= data_in(8487);
     data_out(3588) <= data_in(8491);
     data_out(3589) <= data_in(8493);
     data_out(3590) <= data_in(8495);
     data_out(3591) <= data_in(8500);
     data_out(3592) <= data_in(8501);
     data_out(3593) <= data_in(8504);
     data_out(3594) <= data_in(8505);
     data_out(3595) <= data_in(8506);
     data_out(3596) <= data_in(8509);
     data_out(3597) <= data_in(8512);
     data_out(3598) <= data_in(8516);
     data_out(3599) <= data_in(8519);
     data_out(3600) <= data_in(8523);
     data_out(3601) <= data_in(8525);
     data_out(3602) <= data_in(8527);
     data_out(3603) <= data_in(8530);
     data_out(3604) <= data_in(8531);
     data_out(3605) <= data_in(8533);
     data_out(3606) <= data_in(8535);
     data_out(3607) <= data_in(8536);
     data_out(3608) <= data_in(8539);
     data_out(3609) <= data_in(8540);
     data_out(3610) <= data_in(8543);
     data_out(3611) <= data_in(8544);
     data_out(3612) <= data_in(8546);
     data_out(3613) <= data_in(8547);
     data_out(3614) <= data_in(8548);
     data_out(3615) <= data_in(8554);
     data_out(3616) <= data_in(8555);
     data_out(3617) <= data_in(8557);
     data_out(3618) <= data_in(8562);
     data_out(3619) <= data_in(8569);
     data_out(3620) <= data_in(8570);
     data_out(3621) <= data_in(8573);
     data_out(3622) <= data_in(8576);
     data_out(3623) <= data_in(8579);
     data_out(3624) <= data_in(8580);
     data_out(3625) <= data_in(8581);
     data_out(3626) <= data_in(8585);
     data_out(3627) <= data_in(8592);
     data_out(3628) <= data_in(8593);
     data_out(3629) <= data_in(8595);
     data_out(3630) <= data_in(8596);
     data_out(3631) <= data_in(8597);
     data_out(3632) <= data_in(8601);
     data_out(3633) <= data_in(8603);
     data_out(3634) <= data_in(8606);
     data_out(3635) <= data_in(8607);
     data_out(3636) <= data_in(8612);
     data_out(3637) <= data_in(8622);
     data_out(3638) <= data_in(8623);
     data_out(3639) <= data_in(8626);
     data_out(3640) <= data_in(8628);
     data_out(3641) <= data_in(8633);
     data_out(3642) <= data_in(8636);
     data_out(3643) <= data_in(8638);
     data_out(3644) <= data_in(8639);
     data_out(3645) <= data_in(8642);
     data_out(3646) <= data_in(8647);
     data_out(3647) <= data_in(8648);
     data_out(3648) <= data_in(8655);
     data_out(3649) <= data_in(8656);
     data_out(3650) <= data_in(8660);
     data_out(3651) <= data_in(8661);
     data_out(3652) <= data_in(8663);
     data_out(3653) <= data_in(8668);
     data_out(3654) <= data_in(8669);
     data_out(3655) <= data_in(8671);
     data_out(3656) <= data_in(8675);
     data_out(3657) <= data_in(8676);
     data_out(3658) <= data_in(8680);
     data_out(3659) <= data_in(8683);
     data_out(3660) <= data_in(8686);
     data_out(3661) <= data_in(8687);
     data_out(3662) <= data_in(8688);
     data_out(3663) <= data_in(8690);
     data_out(3664) <= data_in(8692);
     data_out(3665) <= data_in(8693);
     data_out(3666) <= data_in(8694);
     data_out(3667) <= data_in(8696);
     data_out(3668) <= data_in(8697);
     data_out(3669) <= data_in(8700);
     data_out(3670) <= data_in(8703);
     data_out(3671) <= data_in(8705);
     data_out(3672) <= data_in(8711);
     data_out(3673) <= data_in(8712);
     data_out(3674) <= data_in(8717);
     data_out(3675) <= data_in(8718);
     data_out(3676) <= data_in(8723);
     data_out(3677) <= data_in(8725);
     data_out(3678) <= data_in(8726);
     data_out(3679) <= data_in(8727);
     data_out(3680) <= data_in(8730);
     data_out(3681) <= data_in(8731);
     data_out(3682) <= data_in(8734);
     data_out(3683) <= data_in(8735);
     data_out(3684) <= data_in(8741);
     data_out(3685) <= data_in(8743);
     data_out(3686) <= data_in(8745);
     data_out(3687) <= data_in(8746);
     data_out(3688) <= data_in(8750);
     data_out(3689) <= data_in(8751);
     data_out(3690) <= data_in(8758);
     data_out(3691) <= data_in(8763);
     data_out(3692) <= data_in(8764);
     data_out(3693) <= data_in(8769);
     data_out(3694) <= data_in(8772);
     data_out(3695) <= data_in(8774);
     data_out(3696) <= data_in(8780);
     data_out(3697) <= data_in(8781);
     data_out(3698) <= data_in(8783);
     data_out(3699) <= data_in(8784);
     data_out(3700) <= data_in(8785);
     data_out(3701) <= data_in(8787);
     data_out(3702) <= data_in(8788);
     data_out(3703) <= data_in(8792);
     data_out(3704) <= data_in(8795);
     data_out(3705) <= data_in(8797);
     data_out(3706) <= data_in(8799);
     data_out(3707) <= data_in(8801);
     data_out(3708) <= data_in(8802);
     data_out(3709) <= data_in(8803);
     data_out(3710) <= data_in(8804);
     data_out(3711) <= data_in(8805);
     data_out(3712) <= data_in(8806);
     data_out(3713) <= data_in(8808);
     data_out(3714) <= data_in(8809);
     data_out(3715) <= data_in(8810);
     data_out(3716) <= data_in(8814);
     data_out(3717) <= data_in(8817);
     data_out(3718) <= data_in(8818);
     data_out(3719) <= data_in(8819);
     data_out(3720) <= data_in(8820);
     data_out(3721) <= data_in(8822);
     data_out(3722) <= data_in(8825);
     data_out(3723) <= data_in(8826);
     data_out(3724) <= data_in(8827);
     data_out(3725) <= data_in(8828);
     data_out(3726) <= data_in(8832);
     data_out(3727) <= data_in(8833);
     data_out(3728) <= data_in(8836);
     data_out(3729) <= data_in(8837);
     data_out(3730) <= data_in(8838);
     data_out(3731) <= data_in(8846);
     data_out(3732) <= data_in(8847);
     data_out(3733) <= data_in(8848);
     data_out(3734) <= data_in(8849);
     data_out(3735) <= data_in(8851);
     data_out(3736) <= data_in(8852);
     data_out(3737) <= data_in(8853);
     data_out(3738) <= data_in(8854);
     data_out(3739) <= data_in(8855);
     data_out(3740) <= data_in(8858);
     data_out(3741) <= data_in(8859);
     data_out(3742) <= data_in(8862);
     data_out(3743) <= data_in(8864);
     data_out(3744) <= data_in(8869);
     data_out(3745) <= data_in(8876);
     data_out(3746) <= data_in(8878);
     data_out(3747) <= data_in(8880);
     data_out(3748) <= data_in(8883);
     data_out(3749) <= data_in(8884);
     data_out(3750) <= data_in(8885);
     data_out(3751) <= data_in(8886);
     data_out(3752) <= data_in(8887);
     data_out(3753) <= data_in(8890);
     data_out(3754) <= data_in(8892);
     data_out(3755) <= data_in(8893);
     data_out(3756) <= data_in(8899);
     data_out(3757) <= data_in(8901);
     data_out(3758) <= data_in(8903);
     data_out(3759) <= data_in(8904);
     data_out(3760) <= data_in(8907);
     data_out(3761) <= data_in(8908);
     data_out(3762) <= data_in(8909);
     data_out(3763) <= data_in(8913);
     data_out(3764) <= data_in(8914);
     data_out(3765) <= data_in(8918);
     data_out(3766) <= data_in(8922);
     data_out(3767) <= data_in(8923);
     data_out(3768) <= data_in(8926);
     data_out(3769) <= data_in(8928);
     data_out(3770) <= data_in(8929);
     data_out(3771) <= data_in(8933);
     data_out(3772) <= data_in(8934);
     data_out(3773) <= data_in(8937);
     data_out(3774) <= data_in(8938);
     data_out(3775) <= data_in(8939);
     data_out(3776) <= data_in(8948);
     data_out(3777) <= data_in(8951);
     data_out(3778) <= data_in(8968);
     data_out(3779) <= data_in(8970);
     data_out(3780) <= data_in(8977);
     data_out(3781) <= data_in(8979);
     data_out(3782) <= data_in(8980);
     data_out(3783) <= data_in(8981);
     data_out(3784) <= data_in(8982);
     data_out(3785) <= data_in(8991);
     data_out(3786) <= data_in(8992);
     data_out(3787) <= data_in(8995);
     data_out(3788) <= data_in(9005);
     data_out(3789) <= data_in(9006);
     data_out(3790) <= data_in(9012);
     data_out(3791) <= data_in(9014);
     data_out(3792) <= data_in(9017);
     data_out(3793) <= data_in(9020);
     data_out(3794) <= data_in(9029);
     data_out(3795) <= data_in(9030);
     data_out(3796) <= data_in(9034);
     data_out(3797) <= data_in(9038);
     data_out(3798) <= data_in(9043);
     data_out(3799) <= data_in(9044);
     data_out(3800) <= data_in(9045);
     data_out(3801) <= data_in(9046);
     data_out(3802) <= data_in(9054);
     data_out(3803) <= data_in(9060);
     data_out(3804) <= data_in(9061);
     data_out(3805) <= data_in(9062);
     data_out(3806) <= data_in(9064);
     data_out(3807) <= data_in(9066);
     data_out(3808) <= data_in(9067);
     data_out(3809) <= data_in(9070);
     data_out(3810) <= data_in(9076);
     data_out(3811) <= data_in(9078);
     data_out(3812) <= data_in(9079);
     data_out(3813) <= data_in(9080);
     data_out(3814) <= data_in(9082);
     data_out(3815) <= data_in(9085);
     data_out(3816) <= data_in(9087);
     data_out(3817) <= data_in(9090);
     data_out(3818) <= data_in(9095);
     data_out(3819) <= data_in(9097);
     data_out(3820) <= data_in(9101);
     data_out(3821) <= data_in(9102);
     data_out(3822) <= data_in(9103);
     data_out(3823) <= data_in(9107);
     data_out(3824) <= data_in(9108);
     data_out(3825) <= data_in(9109);
     data_out(3826) <= data_in(9114);
     data_out(3827) <= data_in(9116);
     data_out(3828) <= data_in(9118);
     data_out(3829) <= data_in(9119);
     data_out(3830) <= data_in(9121);
     data_out(3831) <= data_in(9123);
     data_out(3832) <= data_in(9124);
     data_out(3833) <= data_in(9126);
     data_out(3834) <= data_in(9131);
     data_out(3835) <= data_in(9138);
     data_out(3836) <= data_in(9140);
     data_out(3837) <= data_in(9142);
     data_out(3838) <= data_in(9143);
     data_out(3839) <= data_in(9148);
     data_out(3840) <= data_in(9155);
     data_out(3841) <= data_in(9157);
     data_out(3842) <= data_in(9162);
     data_out(3843) <= data_in(9164);
     data_out(3844) <= data_in(9166);
     data_out(3845) <= data_in(9168);
     data_out(3846) <= data_in(9170);
     data_out(3847) <= data_in(9175);
     data_out(3848) <= data_in(9176);
     data_out(3849) <= data_in(9178);
     data_out(3850) <= data_in(9180);
     data_out(3851) <= data_in(9181);
     data_out(3852) <= data_in(9182);
     data_out(3853) <= data_in(9184);
     data_out(3854) <= data_in(9188);
     data_out(3855) <= data_in(9193);
     data_out(3856) <= data_in(9194);
     data_out(3857) <= data_in(9196);
     data_out(3858) <= data_in(9197);
     data_out(3859) <= data_in(9198);
     data_out(3860) <= data_in(9199);
     data_out(3861) <= data_in(9201);
     data_out(3862) <= data_in(9204);
     data_out(3863) <= data_in(9205);
     data_out(3864) <= data_in(9206);
     data_out(3865) <= data_in(9207);
     data_out(3866) <= data_in(9208);
     data_out(3867) <= data_in(9212);
     data_out(3868) <= data_in(9213);
     data_out(3869) <= data_in(9217);
     data_out(3870) <= data_in(9218);
     data_out(3871) <= data_in(9219);
     data_out(3872) <= data_in(9221);
     data_out(3873) <= data_in(9222);
     data_out(3874) <= data_in(9223);
     data_out(3875) <= data_in(9231);
     data_out(3876) <= data_in(9234);
     data_out(3877) <= data_in(9235);
     data_out(3878) <= data_in(9236);
     data_out(3879) <= data_in(9238);
     data_out(3880) <= data_in(9244);
     data_out(3881) <= data_in(9249);
     data_out(3882) <= data_in(9252);
     data_out(3883) <= data_in(9253);
     data_out(3884) <= data_in(9255);
     data_out(3885) <= data_in(9263);
     data_out(3886) <= data_in(9266);
     data_out(3887) <= data_in(9267);
     data_out(3888) <= data_in(9269);
     data_out(3889) <= data_in(9271);
     data_out(3890) <= data_in(9273);
     data_out(3891) <= data_in(9274);
     data_out(3892) <= data_in(9276);
     data_out(3893) <= data_in(9277);
     data_out(3894) <= data_in(9278);
     data_out(3895) <= data_in(9279);
     data_out(3896) <= data_in(9281);
     data_out(3897) <= data_in(9282);
     data_out(3898) <= data_in(9284);
     data_out(3899) <= data_in(9286);
     data_out(3900) <= data_in(9287);
     data_out(3901) <= data_in(9289);
     data_out(3902) <= data_in(9292);
     data_out(3903) <= data_in(9293);
     data_out(3904) <= data_in(9298);
     data_out(3905) <= data_in(9302);
     data_out(3906) <= data_in(9307);
     data_out(3907) <= data_in(9309);
     data_out(3908) <= data_in(9315);
     data_out(3909) <= data_in(9316);
     data_out(3910) <= data_in(9318);
     data_out(3911) <= data_in(9319);
     data_out(3912) <= data_in(9323);
     data_out(3913) <= data_in(9324);
     data_out(3914) <= data_in(9325);
     data_out(3915) <= data_in(9327);
     data_out(3916) <= data_in(9328);
     data_out(3917) <= data_in(9330);
     data_out(3918) <= data_in(9331);
     data_out(3919) <= data_in(9333);
     data_out(3920) <= data_in(9335);
     data_out(3921) <= data_in(9337);
     data_out(3922) <= data_in(9338);
     data_out(3923) <= data_in(9339);
     data_out(3924) <= data_in(9341);
     data_out(3925) <= data_in(9347);
     data_out(3926) <= data_in(9348);
     data_out(3927) <= data_in(9349);
     data_out(3928) <= data_in(9350);
     data_out(3929) <= data_in(9351);
     data_out(3930) <= data_in(9352);
     data_out(3931) <= data_in(9354);
     data_out(3932) <= data_in(9355);
     data_out(3933) <= data_in(9356);
     data_out(3934) <= data_in(9360);
     data_out(3935) <= data_in(9361);
     data_out(3936) <= data_in(9367);
     data_out(3937) <= data_in(9369);
     data_out(3938) <= data_in(9370);
     data_out(3939) <= data_in(9374);
     data_out(3940) <= data_in(9375);
     data_out(3941) <= data_in(9379);
     data_out(3942) <= data_in(9382);
     data_out(3943) <= data_in(9383);
     data_out(3944) <= data_in(9387);
     data_out(3945) <= data_in(9388);
     data_out(3946) <= data_in(9391);
     data_out(3947) <= data_in(9401);
     data_out(3948) <= data_in(9402);
     data_out(3949) <= data_in(9403);
     data_out(3950) <= data_in(9405);
     data_out(3951) <= data_in(9406);
     data_out(3952) <= data_in(9407);
     data_out(3953) <= data_in(9409);
     data_out(3954) <= data_in(9410);
     data_out(3955) <= data_in(9411);
     data_out(3956) <= data_in(9412);
     data_out(3957) <= data_in(9415);
     data_out(3958) <= data_in(9416);
     data_out(3959) <= data_in(9417);
     data_out(3960) <= data_in(9419);
     data_out(3961) <= data_in(9424);
     data_out(3962) <= data_in(9425);
     data_out(3963) <= data_in(9429);
     data_out(3964) <= data_in(9431);
     data_out(3965) <= data_in(9432);
     data_out(3966) <= data_in(9433);
     data_out(3967) <= data_in(9435);
     data_out(3968) <= data_in(9438);
     data_out(3969) <= data_in(9441);
     data_out(3970) <= data_in(9445);
     data_out(3971) <= data_in(9448);
     data_out(3972) <= data_in(9451);
     data_out(3973) <= data_in(9452);
     data_out(3974) <= data_in(9456);
     data_out(3975) <= data_in(9458);
     data_out(3976) <= data_in(9460);
     data_out(3977) <= data_in(9462);
     data_out(3978) <= data_in(9466);
     data_out(3979) <= data_in(9470);
     data_out(3980) <= data_in(9478);
     data_out(3981) <= data_in(9483);
     data_out(3982) <= data_in(9485);
     data_out(3983) <= data_in(9486);
     data_out(3984) <= data_in(9487);
     data_out(3985) <= data_in(9489);
     data_out(3986) <= data_in(9490);
     data_out(3987) <= data_in(9494);
     data_out(3988) <= data_in(9495);
     data_out(3989) <= data_in(9496);
     data_out(3990) <= data_in(9500);
     data_out(3991) <= data_in(9502);
     data_out(3992) <= data_in(9503);
     data_out(3993) <= data_in(9509);
     data_out(3994) <= data_in(9510);
     data_out(3995) <= data_in(9511);
     data_out(3996) <= data_in(9512);
     data_out(3997) <= data_in(9513);
     data_out(3998) <= data_in(9516);
     data_out(3999) <= data_in(9520);
     data_out(4000) <= data_in(9521);
     data_out(4001) <= data_in(9524);
     data_out(4002) <= data_in(9528);
     data_out(4003) <= data_in(9529);
     data_out(4004) <= data_in(9533);
     data_out(4005) <= data_in(9536);
     data_out(4006) <= data_in(9542);
     data_out(4007) <= data_in(9544);
     data_out(4008) <= data_in(9550);
     data_out(4009) <= data_in(9551);
     data_out(4010) <= data_in(9555);
     data_out(4011) <= data_in(9558);
     data_out(4012) <= data_in(9560);
     data_out(4013) <= data_in(9563);
     data_out(4014) <= data_in(9565);
     data_out(4015) <= data_in(9567);
     data_out(4016) <= data_in(9570);
     data_out(4017) <= data_in(9575);
     data_out(4018) <= data_in(9578);
     data_out(4019) <= data_in(9579);
     data_out(4020) <= data_in(9583);
     data_out(4021) <= data_in(9585);
     data_out(4022) <= data_in(9587);
     data_out(4023) <= data_in(9591);
     data_out(4024) <= data_in(9593);
     data_out(4025) <= data_in(9594);
     data_out(4026) <= data_in(9595);
     data_out(4027) <= data_in(9600);
     data_out(4028) <= data_in(9602);
     data_out(4029) <= data_in(9603);
     data_out(4030) <= data_in(9604);
     data_out(4031) <= data_in(9607);
     data_out(4032) <= data_in(9609);
     data_out(4033) <= data_in(9616);
     data_out(4034) <= data_in(9624);
     data_out(4035) <= data_in(9631);
     data_out(4036) <= data_in(9632);
     data_out(4037) <= data_in(9635);
     data_out(4038) <= data_in(9636);
     data_out(4039) <= data_in(9640);
     data_out(4040) <= data_in(9644);
     data_out(4041) <= data_in(9647);
     data_out(4042) <= data_in(9650);
     data_out(4043) <= data_in(9653);
     data_out(4044) <= data_in(9657);
     data_out(4045) <= data_in(9663);
     data_out(4046) <= data_in(9667);
     data_out(4047) <= data_in(9672);
     data_out(4048) <= data_in(9673);
     data_out(4049) <= data_in(9675);
     data_out(4050) <= data_in(9679);
     data_out(4051) <= data_in(9681);
     data_out(4052) <= data_in(9682);
     data_out(4053) <= data_in(9685);
     data_out(4054) <= data_in(9686);
     data_out(4055) <= data_in(9688);
     data_out(4056) <= data_in(9691);
     data_out(4057) <= data_in(9693);
     data_out(4058) <= data_in(9696);
     data_out(4059) <= data_in(9698);
     data_out(4060) <= data_in(9701);
     data_out(4061) <= data_in(9703);
     data_out(4062) <= data_in(9709);
     data_out(4063) <= data_in(9710);
     data_out(4064) <= data_in(9711);
     data_out(4065) <= data_in(9713);
     data_out(4066) <= data_in(9714);
     data_out(4067) <= data_in(9716);
     data_out(4068) <= data_in(9718);
     data_out(4069) <= data_in(9719);
     data_out(4070) <= data_in(9722);
     data_out(4071) <= data_in(9727);
     data_out(4072) <= data_in(9728);
     data_out(4073) <= data_in(9740);
     data_out(4074) <= data_in(9742);
     data_out(4075) <= data_in(9745);
     data_out(4076) <= data_in(9746);
     data_out(4077) <= data_in(9755);
     data_out(4078) <= data_in(9759);
     data_out(4079) <= data_in(9762);
     data_out(4080) <= data_in(9766);
     data_out(4081) <= data_in(9767);
     data_out(4082) <= data_in(9769);
     data_out(4083) <= data_in(9773);
     data_out(4084) <= data_in(9774);
     data_out(4085) <= data_in(9780);
     data_out(4086) <= data_in(9781);
     data_out(4087) <= data_in(9783);
     data_out(4088) <= data_in(9784);
     data_out(4089) <= data_in(9786);
     data_out(4090) <= data_in(9787);
     data_out(4091) <= data_in(9797);
     data_out(4092) <= data_in(9799);
     data_out(4093) <= data_in(9805);
     data_out(4094) <= data_in(9809);
     data_out(4095) <= data_in(9810);
     data_out(4096) <= data_in(9811);
     data_out(4097) <= data_in(9813);
     data_out(4098) <= data_in(9814);
     data_out(4099) <= data_in(9818);
     data_out(4100) <= data_in(9821);
     data_out(4101) <= data_in(9824);
     data_out(4102) <= data_in(9825);
     data_out(4103) <= data_in(9828);
     data_out(4104) <= data_in(9829);
     data_out(4105) <= data_in(9832);
     data_out(4106) <= data_in(9835);
     data_out(4107) <= data_in(9838);
     data_out(4108) <= data_in(9839);
     data_out(4109) <= data_in(9842);
     data_out(4110) <= data_in(9847);
     data_out(4111) <= data_in(9851);
     data_out(4112) <= data_in(9857);
     data_out(4113) <= data_in(9861);
     data_out(4114) <= data_in(9863);
     data_out(4115) <= data_in(9871);
     data_out(4116) <= data_in(9875);
     data_out(4117) <= data_in(9880);
     data_out(4118) <= data_in(9881);
     data_out(4119) <= data_in(9882);
     data_out(4120) <= data_in(9884);
     data_out(4121) <= data_in(9885);
     data_out(4122) <= data_in(9887);
     data_out(4123) <= data_in(9888);
     data_out(4124) <= data_in(9893);
     data_out(4125) <= data_in(9897);
     data_out(4126) <= data_in(9899);
     data_out(4127) <= data_in(9900);
     data_out(4128) <= data_in(9902);
     data_out(4129) <= data_in(9904);
     data_out(4130) <= data_in(9908);
     data_out(4131) <= data_in(9909);
     data_out(4132) <= data_in(9911);
     data_out(4133) <= data_in(9913);
     data_out(4134) <= data_in(9914);
     data_out(4135) <= data_in(9920);
     data_out(4136) <= data_in(9923);
     data_out(4137) <= data_in(9925);
     data_out(4138) <= data_in(9926);
     data_out(4139) <= data_in(9932);
     data_out(4140) <= data_in(9935);
     data_out(4141) <= data_in(9937);
     data_out(4142) <= data_in(9938);
     data_out(4143) <= data_in(9941);
     data_out(4144) <= data_in(9942);
     data_out(4145) <= data_in(9943);
     data_out(4146) <= data_in(9944);
     data_out(4147) <= data_in(9947);
     data_out(4148) <= data_in(9949);
     data_out(4149) <= data_in(9953);
     data_out(4150) <= data_in(9955);
     data_out(4151) <= data_in(9959);
     data_out(4152) <= data_in(9960);
     data_out(4153) <= data_in(9961);
     data_out(4154) <= data_in(9962);
     data_out(4155) <= data_in(9965);
     data_out(4156) <= data_in(9966);
     data_out(4157) <= data_in(9968);
     data_out(4158) <= data_in(9970);
     data_out(4159) <= data_in(9972);
     data_out(4160) <= data_in(9973);
     data_out(4161) <= data_in(9975);
     data_out(4162) <= data_in(9979);
     data_out(4163) <= data_in(9980);
     data_out(4164) <= data_in(9981);
     data_out(4165) <= data_in(9983);
     data_out(4166) <= data_in(9986);
     data_out(4167) <= data_in(9987);
     data_out(4168) <= data_in(9988);
     data_out(4169) <= data_in(9989);
     data_out(4170) <= data_in(9990);
     data_out(4171) <= data_in(9991);
     data_out(4172) <= data_in(9996);
     data_out(4173) <= data_in(9999);
     data_out(4174) <= data_in(10000);
     data_out(4175) <= data_in(10003);
     data_out(4176) <= data_in(10007);
     data_out(4177) <= data_in(10013);
     data_out(4178) <= data_in(10019);
     data_out(4179) <= data_in(10025);
     data_out(4180) <= data_in(10027);
     data_out(4181) <= data_in(10028);
     data_out(4182) <= data_in(10029);
     data_out(4183) <= data_in(10031);
     data_out(4184) <= data_in(10032);
     data_out(4185) <= data_in(10038);
     data_out(4186) <= data_in(10040);
     data_out(4187) <= data_in(10042);
     data_out(4188) <= data_in(10047);
     data_out(4189) <= data_in(10049);
     data_out(4190) <= data_in(10051);
     data_out(4191) <= data_in(10052);
     data_out(4192) <= data_in(10053);
     data_out(4193) <= data_in(10060);
     data_out(4194) <= data_in(10061);
     data_out(4195) <= data_in(10062);
     data_out(4196) <= data_in(10066);
     data_out(4197) <= data_in(10070);
     data_out(4198) <= data_in(10072);
     data_out(4199) <= data_in(10073);
     data_out(4200) <= data_in(10074);
     data_out(4201) <= data_in(10075);
     data_out(4202) <= data_in(10078);
     data_out(4203) <= data_in(10079);
     data_out(4204) <= data_in(10080);
     data_out(4205) <= data_in(10081);
     data_out(4206) <= data_in(10083);
     data_out(4207) <= data_in(10084);
     data_out(4208) <= data_in(10086);
     data_out(4209) <= data_in(10093);
     data_out(4210) <= data_in(10094);
     data_out(4211) <= data_in(10095);
     data_out(4212) <= data_in(10096);
     data_out(4213) <= data_in(10098);
     data_out(4214) <= data_in(10102);
     data_out(4215) <= data_in(10103);
     data_out(4216) <= data_in(10106);
     data_out(4217) <= data_in(10112);
     data_out(4218) <= data_in(10113);
     data_out(4219) <= data_in(10115);
     data_out(4220) <= data_in(10118);
     data_out(4221) <= data_in(10119);
     data_out(4222) <= data_in(10120);
     data_out(4223) <= data_in(10122);
     data_out(4224) <= data_in(10126);
     data_out(4225) <= data_in(10131);
     data_out(4226) <= data_in(10132);
     data_out(4227) <= data_in(10138);
     data_out(4228) <= data_in(10139);
     data_out(4229) <= data_in(10141);
     data_out(4230) <= data_in(10142);
     data_out(4231) <= data_in(10145);
     data_out(4232) <= data_in(10151);
     data_out(4233) <= data_in(10153);
     data_out(4234) <= data_in(10164);
     data_out(4235) <= data_in(10165);
     data_out(4236) <= data_in(10171);
     data_out(4237) <= data_in(10177);
     data_out(4238) <= data_in(10181);
     data_out(4239) <= data_in(10182);
     data_out(4240) <= data_in(10186);
     data_out(4241) <= data_in(10187);
     data_out(4242) <= data_in(10188);
     data_out(4243) <= data_in(10198);
     data_out(4244) <= data_in(10199);
     data_out(4245) <= data_in(10200);
     data_out(4246) <= data_in(10203);
     data_out(4247) <= data_in(10204);
     data_out(4248) <= data_in(10205);
     data_out(4249) <= data_in(10206);
     data_out(4250) <= data_in(10207);
     data_out(4251) <= data_in(10209);
     data_out(4252) <= data_in(10210);
     data_out(4253) <= data_in(10216);
     data_out(4254) <= data_in(10219);
     data_out(4255) <= data_in(10225);
     data_out(4256) <= data_in(10228);
     data_out(4257) <= data_in(10229);
     data_out(4258) <= data_in(10230);
     data_out(4259) <= data_in(10235);
     data_out(4260) <= data_in(328);
     data_out(4261) <= data_in(368);
     data_out(4262) <= data_in(466);
     data_out(4263) <= data_in(481);
     data_out(4264) <= data_in(716);
     data_out(4265) <= data_in(772);
     data_out(4266) <= data_in(774);
     data_out(4267) <= data_in(991);
     data_out(4268) <= data_in(1066);
     data_out(4269) <= data_in(1432);
     data_out(4270) <= data_in(1629);
     data_out(4271) <= data_in(1734);
     data_out(4272) <= data_in(1794);
     data_out(4273) <= data_in(1862);
     data_out(4274) <= data_in(1867);
     data_out(4275) <= data_in(1975);
     data_out(4276) <= data_in(2142);
     data_out(4277) <= data_in(2274);
     data_out(4278) <= data_in(2666);
     data_out(4279) <= data_in(2830);
     data_out(4280) <= data_in(2925);
     data_out(4281) <= data_in(2965);
     data_out(4282) <= data_in(3060);
     data_out(4283) <= data_in(3091);
     data_out(4284) <= data_in(3093);
     data_out(4285) <= data_in(3395);
     data_out(4286) <= data_in(3422);
     data_out(4287) <= data_in(3646);
     data_out(4288) <= data_in(4257);
     data_out(4289) <= data_in(4409);
     data_out(4290) <= data_in(4519);
     data_out(4291) <= data_in(4566);
     data_out(4292) <= data_in(4914);
     data_out(4293) <= data_in(4917);
     data_out(4294) <= data_in(5024);
     data_out(4295) <= data_in(5177);
     data_out(4296) <= data_in(5254);
     data_out(4297) <= data_in(5369);
     data_out(4298) <= data_in(5714);
     data_out(4299) <= data_in(6006);
     data_out(4300) <= data_in(6275);
     data_out(4301) <= data_in(6328);
     data_out(4302) <= data_in(6337);
     data_out(4303) <= data_in(6354);
     data_out(4304) <= data_in(6389);
     data_out(4305) <= data_in(6605);
     data_out(4306) <= data_in(6652);
     data_out(4307) <= data_in(7152);
     data_out(4308) <= data_in(7169);
     data_out(4309) <= data_in(7177);
     data_out(4310) <= data_in(7324);
     data_out(4311) <= data_in(7381);
     data_out(4312) <= data_in(7509);
     data_out(4313) <= data_in(7840);
     data_out(4314) <= data_in(8116);
     data_out(4315) <= data_in(8171);
     data_out(4316) <= data_in(8303);
     data_out(4317) <= data_in(8325);
     data_out(4318) <= data_in(8348);
     data_out(4319) <= data_in(8481);
     data_out(4320) <= data_in(8600);
     data_out(4321) <= data_in(8605);
     data_out(4322) <= data_in(8714);
     data_out(4323) <= data_in(8842);
     data_out(4324) <= data_in(8872);
     data_out(4325) <= data_in(9077);
     data_out(4326) <= data_in(9258);
     data_out(4327) <= data_in(9605);
     data_out(4328) <= data_in(9735);
     data_out(4329) <= data_in(9739);
     data_out(4330) <= data_in(9872);
     data_out(4331) <= data_in(9889);
     data_out(4332) <= data_in(9945);
     data_out(4333) <= data_in(10021);
     data_out(4334) <= data_in(10023);
     data_out(4335) <= data_in(10039);
     data_out(4336) <= data_in(10065);
     data_out(4337) <= data_in(10218);
     data_out(4338) <= data_in(288);
     data_out(4339) <= data_in(662);
     data_out(4340) <= data_in(999);
     data_out(4341) <= data_in(1085);
     data_out(4342) <= data_in(1132);
     data_out(4343) <= data_in(1694);
     data_out(4344) <= data_in(1796);
     data_out(4345) <= data_in(1951);
     data_out(4346) <= data_in(2138);
     data_out(4347) <= data_in(2278);
     data_out(4348) <= data_in(2587);
     data_out(4349) <= data_in(2671);
     data_out(4350) <= data_in(2939);
     data_out(4351) <= data_in(3375);
     data_out(4352) <= data_in(3400);
     data_out(4353) <= data_in(3662);
     data_out(4354) <= data_in(3720);
     data_out(4355) <= data_in(3919);
     data_out(4356) <= data_in(3936);
     data_out(4357) <= data_in(3954);
     data_out(4358) <= data_in(3960);
     data_out(4359) <= data_in(4044);
     data_out(4360) <= data_in(4048);
     data_out(4361) <= data_in(4287);
     data_out(4362) <= data_in(4312);
     data_out(4363) <= data_in(4523);
     data_out(4364) <= data_in(4605);
     data_out(4365) <= data_in(4647);
     data_out(4366) <= data_in(4825);
     data_out(4367) <= data_in(4919);
     data_out(4368) <= data_in(5165);
     data_out(4369) <= data_in(5451);
     data_out(4370) <= data_in(5561);
     data_out(4371) <= data_in(5795);
     data_out(4372) <= data_in(5934);
     data_out(4373) <= data_in(6266);
     data_out(4374) <= data_in(6278);
     data_out(4375) <= data_in(6362);
     data_out(4376) <= data_in(6438);
     data_out(4377) <= data_in(6472);
     data_out(4378) <= data_in(6626);
     data_out(4379) <= data_in(7123);
     data_out(4380) <= data_in(7890);
     data_out(4381) <= data_in(8090);
     data_out(4382) <= data_in(8434);
     data_out(4383) <= data_in(8610);
     data_out(4384) <= data_in(9133);
     data_out(4385) <= data_in(9306);
     data_out(4386) <= data_in(9427);
     data_out(4387) <= data_in(9756);
     data_out(4388) <= data_in(10172);
     data_out(4389) <= data_in(10180);
     data_out(4390) <= data_in(240);
     data_out(4391) <= data_in(438);
     data_out(4392) <= data_in(604);
     data_out(4393) <= data_in(952);
     data_out(4394) <= data_in(1133);
     data_out(4395) <= data_in(1697);
     data_out(4396) <= data_in(2004);
     data_out(4397) <= data_in(2125);
     data_out(4398) <= data_in(2212);
     data_out(4399) <= data_in(2280);
     data_out(4400) <= data_in(2368);
     data_out(4401) <= data_in(2499);
     data_out(4402) <= data_in(2711);
     data_out(4403) <= data_in(2810);
     data_out(4404) <= data_in(2987);
     data_out(4405) <= data_in(3278);
     data_out(4406) <= data_in(3329);
     data_out(4407) <= data_in(3391);
     data_out(4408) <= data_in(3535);
     data_out(4409) <= data_in(3601);
     data_out(4410) <= data_in(3647);
     data_out(4411) <= data_in(3652);
     data_out(4412) <= data_in(3691);
     data_out(4413) <= data_in(3753);
     data_out(4414) <= data_in(4388);
     data_out(4415) <= data_in(4489);
     data_out(4416) <= data_in(4511);
     data_out(4417) <= data_in(4561);
     data_out(4418) <= data_in(4590);
     data_out(4419) <= data_in(4868);
     data_out(4420) <= data_in(4928);
     data_out(4421) <= data_in(5295);
     data_out(4422) <= data_in(5469);
     data_out(4423) <= data_in(5538);
     data_out(4424) <= data_in(5673);
     data_out(4425) <= data_in(5741);
     data_out(4426) <= data_in(5838);
     data_out(4427) <= data_in(6002);
     data_out(4428) <= data_in(6005);
     data_out(4429) <= data_in(6049);
     data_out(4430) <= data_in(6171);
     data_out(4431) <= data_in(6282);
     data_out(4432) <= data_in(6833);
     data_out(4433) <= data_in(7057);
     data_out(4434) <= data_in(7126);
     data_out(4435) <= data_in(7218);
     data_out(4436) <= data_in(7336);
     data_out(4437) <= data_in(7373);
     data_out(4438) <= data_in(7493);
     data_out(4439) <= data_in(7947);
     data_out(4440) <= data_in(8173);
     data_out(4441) <= data_in(8193);
     data_out(4442) <= data_in(8197);
     data_out(4443) <= data_in(8237);
     data_out(4444) <= data_in(8662);
     data_out(4445) <= data_in(8944);
     data_out(4446) <= data_in(9001);
     data_out(4447) <= data_in(9147);
     data_out(4448) <= data_in(9668);
     data_out(4449) <= data_in(9748);
     data_out(4450) <= data_in(9982);
     data_out(4451) <= data_in(558);
     data_out(4452) <= data_in(622);
     data_out(4453) <= data_in(654);
     data_out(4454) <= data_in(663);
     data_out(4455) <= data_in(747);
     data_out(4456) <= data_in(854);
     data_out(4457) <= data_in(918);
     data_out(4458) <= data_in(1025);
     data_out(4459) <= data_in(1107);
     data_out(4460) <= data_in(1205);
     data_out(4461) <= data_in(1339);
     data_out(4462) <= data_in(1374);
     data_out(4463) <= data_in(1436);
     data_out(4464) <= data_in(1805);
     data_out(4465) <= data_in(2214);
     data_out(4466) <= data_in(2331);
     data_out(4467) <= data_in(2375);
     data_out(4468) <= data_in(2752);
     data_out(4469) <= data_in(3027);
     data_out(4470) <= data_in(3106);
     data_out(4471) <= data_in(3374);
     data_out(4472) <= data_in(3545);
     data_out(4473) <= data_in(3611);
     data_out(4474) <= data_in(3758);
     data_out(4475) <= data_in(4393);
     data_out(4476) <= data_in(5053);
     data_out(4477) <= data_in(5273);
     data_out(4478) <= data_in(5408);
     data_out(4479) <= data_in(5841);
     data_out(4480) <= data_in(6077);
     data_out(4481) <= data_in(6107);
     data_out(4482) <= data_in(6305);
     data_out(4483) <= data_in(6734);
     data_out(4484) <= data_in(6752);
     data_out(4485) <= data_in(7709);
     data_out(4486) <= data_in(7967);
     data_out(4487) <= data_in(8427);
     data_out(4488) <= data_in(8537);
     data_out(4489) <= data_in(8728);
     data_out(4490) <= data_in(8942);
     data_out(4491) <= data_in(8949);
     data_out(4492) <= data_in(9841);
     data_out(4493) <= data_in(9906);
     data_out(4494) <= data_in(10104);
     data_out(4495) <= data_in(10173);
     data_out(4496) <= data_in(350);
     data_out(4497) <= data_in(352);
     data_out(4498) <= data_in(569);
     data_out(4499) <= data_in(873);
     data_out(4500) <= data_in(934);
     data_out(4501) <= data_in(1529);
     data_out(4502) <= data_in(1558);
     data_out(4503) <= data_in(1616);
     data_out(4504) <= data_in(1666);
     data_out(4505) <= data_in(1837);
     data_out(4506) <= data_in(1860);
     data_out(4507) <= data_in(1873);
     data_out(4508) <= data_in(2361);
     data_out(4509) <= data_in(2588);
     data_out(4510) <= data_in(2593);
     data_out(4511) <= data_in(2657);
     data_out(4512) <= data_in(2880);
     data_out(4513) <= data_in(2900);
     data_out(4514) <= data_in(3405);
     data_out(4515) <= data_in(3438);
     data_out(4516) <= data_in(3579);
     data_out(4517) <= data_in(3749);
     data_out(4518) <= data_in(4361);
     data_out(4519) <= data_in(4540);
     data_out(4520) <= data_in(4691);
     data_out(4521) <= data_in(4816);
     data_out(4522) <= data_in(4905);
     data_out(4523) <= data_in(5083);
     data_out(4524) <= data_in(5185);
     data_out(4525) <= data_in(5323);
     data_out(4526) <= data_in(5604);
     data_out(4527) <= data_in(5719);
     data_out(4528) <= data_in(5761);
     data_out(4529) <= data_in(5794);
     data_out(4530) <= data_in(5960);
     data_out(4531) <= data_in(6452);
     data_out(4532) <= data_in(6736);
     data_out(4533) <= data_in(7374);
     data_out(4534) <= data_in(7392);
     data_out(4535) <= data_in(7669);
     data_out(4536) <= data_in(7723);
     data_out(4537) <= data_in(7832);
     data_out(4538) <= data_in(7938);
     data_out(4539) <= data_in(7972);
     data_out(4540) <= data_in(8100);
     data_out(4541) <= data_in(8105);
     data_out(4542) <= data_in(8286);
     data_out(4543) <= data_in(8398);
     data_out(4544) <= data_in(8964);
     data_out(4545) <= data_in(9240);
     data_out(4546) <= data_in(9480);
     data_out(4547) <= data_in(9771);
     data_out(4548) <= data_in(9791);
     data_out(4549) <= data_in(9860);
     data_out(4550) <= data_in(9930);
     data_out(4551) <= data_in(10152);
     data_out(4552) <= data_in(10214);
     data_out(4553) <= data_in(241);
     data_out(4554) <= data_in(242);
     data_out(4555) <= data_in(244);
     data_out(4556) <= data_in(245);
     data_out(4557) <= data_in(247);
     data_out(4558) <= data_in(253);
     data_out(4559) <= data_in(254);
     data_out(4560) <= data_in(255);
     data_out(4561) <= data_in(256);
     data_out(4562) <= data_in(263);
     data_out(4563) <= data_in(264);
     data_out(4564) <= data_in(267);
     data_out(4565) <= data_in(269);
     data_out(4566) <= data_in(270);
     data_out(4567) <= data_in(272);
     data_out(4568) <= data_in(273);
     data_out(4569) <= data_in(274);
     data_out(4570) <= data_in(275);
     data_out(4571) <= data_in(276);
     data_out(4572) <= data_in(278);
     data_out(4573) <= data_in(285);
     data_out(4574) <= data_in(287);
     data_out(4575) <= data_in(289);
     data_out(4576) <= data_in(293);
     data_out(4577) <= data_in(296);
     data_out(4578) <= data_in(297);
     data_out(4579) <= data_in(298);
     data_out(4580) <= data_in(300);
     data_out(4581) <= data_in(301);
     data_out(4582) <= data_in(302);
     data_out(4583) <= data_in(303);
     data_out(4584) <= data_in(306);
     data_out(4585) <= data_in(308);
     data_out(4586) <= data_in(309);
     data_out(4587) <= data_in(310);
     data_out(4588) <= data_in(312);
     data_out(4589) <= data_in(315);
     data_out(4590) <= data_in(316);
     data_out(4591) <= data_in(317);
     data_out(4592) <= data_in(321);
     data_out(4593) <= data_in(333);
     data_out(4594) <= data_in(335);
     data_out(4595) <= data_in(337);
     data_out(4596) <= data_in(338);
     data_out(4597) <= data_in(339);
     data_out(4598) <= data_in(340);
     data_out(4599) <= data_in(341);
     data_out(4600) <= data_in(342);
     data_out(4601) <= data_in(346);
     data_out(4602) <= data_in(348);
     data_out(4603) <= data_in(351);
     data_out(4604) <= data_in(357);
     data_out(4605) <= data_in(358);
     data_out(4606) <= data_in(363);
     data_out(4607) <= data_in(365);
     data_out(4608) <= data_in(366);
     data_out(4609) <= data_in(373);
     data_out(4610) <= data_in(374);
     data_out(4611) <= data_in(375);
     data_out(4612) <= data_in(376);
     data_out(4613) <= data_in(377);
     data_out(4614) <= data_in(380);
     data_out(4615) <= data_in(382);
     data_out(4616) <= data_in(383);
     data_out(4617) <= data_in(385);
     data_out(4618) <= data_in(386);
     data_out(4619) <= data_in(390);
     data_out(4620) <= data_in(392);
     data_out(4621) <= data_in(395);
     data_out(4622) <= data_in(397);
     data_out(4623) <= data_in(398);
     data_out(4624) <= data_in(401);
     data_out(4625) <= data_in(402);
     data_out(4626) <= data_in(403);
     data_out(4627) <= data_in(404);
     data_out(4628) <= data_in(407);
     data_out(4629) <= data_in(410);
     data_out(4630) <= data_in(415);
     data_out(4631) <= data_in(416);
     data_out(4632) <= data_in(418);
     data_out(4633) <= data_in(421);
     data_out(4634) <= data_in(422);
     data_out(4635) <= data_in(425);
     data_out(4636) <= data_in(427);
     data_out(4637) <= data_in(430);
     data_out(4638) <= data_in(431);
     data_out(4639) <= data_in(436);
     data_out(4640) <= data_in(443);
     data_out(4641) <= data_in(448);
     data_out(4642) <= data_in(451);
     data_out(4643) <= data_in(453);
     data_out(4644) <= data_in(454);
     data_out(4645) <= data_in(455);
     data_out(4646) <= data_in(457);
     data_out(4647) <= data_in(460);
     data_out(4648) <= data_in(464);
     data_out(4649) <= data_in(472);
     data_out(4650) <= data_in(475);
     data_out(4651) <= data_in(476);
     data_out(4652) <= data_in(479);
     data_out(4653) <= data_in(482);
     data_out(4654) <= data_in(484);
     data_out(4655) <= data_in(490);
     data_out(4656) <= data_in(491);
     data_out(4657) <= data_in(494);
     data_out(4658) <= data_in(496);
     data_out(4659) <= data_in(497);
     data_out(4660) <= data_in(498);
     data_out(4661) <= data_in(499);
     data_out(4662) <= data_in(501);
     data_out(4663) <= data_in(503);
     data_out(4664) <= data_in(506);
     data_out(4665) <= data_in(508);
     data_out(4666) <= data_in(512);
     data_out(4667) <= data_in(515);
     data_out(4668) <= data_in(517);
     data_out(4669) <= data_in(518);
     data_out(4670) <= data_in(519);
     data_out(4671) <= data_in(523);
     data_out(4672) <= data_in(525);
     data_out(4673) <= data_in(526);
     data_out(4674) <= data_in(527);
     data_out(4675) <= data_in(529);
     data_out(4676) <= data_in(530);
     data_out(4677) <= data_in(531);
     data_out(4678) <= data_in(532);
     data_out(4679) <= data_in(536);
     data_out(4680) <= data_in(540);
     data_out(4681) <= data_in(543);
     data_out(4682) <= data_in(550);
     data_out(4683) <= data_in(552);
     data_out(4684) <= data_in(557);
     data_out(4685) <= data_in(561);
     data_out(4686) <= data_in(564);
     data_out(4687) <= data_in(565);
     data_out(4688) <= data_in(573);
     data_out(4689) <= data_in(575);
     data_out(4690) <= data_in(581);
     data_out(4691) <= data_in(584);
     data_out(4692) <= data_in(587);
     data_out(4693) <= data_in(592);
     data_out(4694) <= data_in(597);
     data_out(4695) <= data_in(610);
     data_out(4696) <= data_in(611);
     data_out(4697) <= data_in(616);
     data_out(4698) <= data_in(617);
     data_out(4699) <= data_in(618);
     data_out(4700) <= data_in(625);
     data_out(4701) <= data_in(627);
     data_out(4702) <= data_in(628);
     data_out(4703) <= data_in(634);
     data_out(4704) <= data_in(635);
     data_out(4705) <= data_in(638);
     data_out(4706) <= data_in(640);
     data_out(4707) <= data_in(641);
     data_out(4708) <= data_in(644);
     data_out(4709) <= data_in(645);
     data_out(4710) <= data_in(646);
     data_out(4711) <= data_in(650);
     data_out(4712) <= data_in(651);
     data_out(4713) <= data_in(652);
     data_out(4714) <= data_in(655);
     data_out(4715) <= data_in(664);
     data_out(4716) <= data_in(665);
     data_out(4717) <= data_in(666);
     data_out(4718) <= data_in(667);
     data_out(4719) <= data_in(675);
     data_out(4720) <= data_in(680);
     data_out(4721) <= data_in(684);
     data_out(4722) <= data_in(686);
     data_out(4723) <= data_in(688);
     data_out(4724) <= data_in(689);
     data_out(4725) <= data_in(690);
     data_out(4726) <= data_in(691);
     data_out(4727) <= data_in(693);
     data_out(4728) <= data_in(696);
     data_out(4729) <= data_in(701);
     data_out(4730) <= data_in(703);
     data_out(4731) <= data_in(704);
     data_out(4732) <= data_in(705);
     data_out(4733) <= data_in(707);
     data_out(4734) <= data_in(709);
     data_out(4735) <= data_in(710);
     data_out(4736) <= data_in(712);
     data_out(4737) <= data_in(717);
     data_out(4738) <= data_in(718);
     data_out(4739) <= data_in(720);
     data_out(4740) <= data_in(721);
     data_out(4741) <= data_in(723);
     data_out(4742) <= data_in(724);
     data_out(4743) <= data_in(729);
     data_out(4744) <= data_in(730);
     data_out(4745) <= data_in(731);
     data_out(4746) <= data_in(733);
     data_out(4747) <= data_in(740);
     data_out(4748) <= data_in(742);
     data_out(4749) <= data_in(745);
     data_out(4750) <= data_in(746);
     data_out(4751) <= data_in(750);
     data_out(4752) <= data_in(751);
     data_out(4753) <= data_in(756);
     data_out(4754) <= data_in(765);
     data_out(4755) <= data_in(766);
     data_out(4756) <= data_in(767);
     data_out(4757) <= data_in(775);
     data_out(4758) <= data_in(777);
     data_out(4759) <= data_in(779);
     data_out(4760) <= data_in(780);
     data_out(4761) <= data_in(787);
     data_out(4762) <= data_in(790);
     data_out(4763) <= data_in(792);
     data_out(4764) <= data_in(793);
     data_out(4765) <= data_in(794);
     data_out(4766) <= data_in(795);
     data_out(4767) <= data_in(796);
     data_out(4768) <= data_in(800);
     data_out(4769) <= data_in(802);
     data_out(4770) <= data_in(807);
     data_out(4771) <= data_in(809);
     data_out(4772) <= data_in(811);
     data_out(4773) <= data_in(812);
     data_out(4774) <= data_in(813);
     data_out(4775) <= data_in(816);
     data_out(4776) <= data_in(819);
     data_out(4777) <= data_in(822);
     data_out(4778) <= data_in(824);
     data_out(4779) <= data_in(826);
     data_out(4780) <= data_in(827);
     data_out(4781) <= data_in(828);
     data_out(4782) <= data_in(832);
     data_out(4783) <= data_in(833);
     data_out(4784) <= data_in(834);
     data_out(4785) <= data_in(844);
     data_out(4786) <= data_in(846);
     data_out(4787) <= data_in(847);
     data_out(4788) <= data_in(850);
     data_out(4789) <= data_in(851);
     data_out(4790) <= data_in(852);
     data_out(4791) <= data_in(855);
     data_out(4792) <= data_in(856);
     data_out(4793) <= data_in(857);
     data_out(4794) <= data_in(859);
     data_out(4795) <= data_in(860);
     data_out(4796) <= data_in(861);
     data_out(4797) <= data_in(867);
     data_out(4798) <= data_in(869);
     data_out(4799) <= data_in(871);
     data_out(4800) <= data_in(875);
     data_out(4801) <= data_in(877);
     data_out(4802) <= data_in(880);
     data_out(4803) <= data_in(883);
     data_out(4804) <= data_in(887);
     data_out(4805) <= data_in(890);
     data_out(4806) <= data_in(891);
     data_out(4807) <= data_in(892);
     data_out(4808) <= data_in(896);
     data_out(4809) <= data_in(901);
     data_out(4810) <= data_in(902);
     data_out(4811) <= data_in(903);
     data_out(4812) <= data_in(904);
     data_out(4813) <= data_in(905);
     data_out(4814) <= data_in(906);
     data_out(4815) <= data_in(907);
     data_out(4816) <= data_in(908);
     data_out(4817) <= data_in(909);
     data_out(4818) <= data_in(911);
     data_out(4819) <= data_in(912);
     data_out(4820) <= data_in(915);
     data_out(4821) <= data_in(917);
     data_out(4822) <= data_in(922);
     data_out(4823) <= data_in(933);
     data_out(4824) <= data_in(937);
     data_out(4825) <= data_in(941);
     data_out(4826) <= data_in(944);
     data_out(4827) <= data_in(945);
     data_out(4828) <= data_in(947);
     data_out(4829) <= data_in(951);
     data_out(4830) <= data_in(954);
     data_out(4831) <= data_in(955);
     data_out(4832) <= data_in(956);
     data_out(4833) <= data_in(957);
     data_out(4834) <= data_in(958);
     data_out(4835) <= data_in(959);
     data_out(4836) <= data_in(962);
     data_out(4837) <= data_in(974);
     data_out(4838) <= data_in(976);
     data_out(4839) <= data_in(978);
     data_out(4840) <= data_in(981);
     data_out(4841) <= data_in(987);
     data_out(4842) <= data_in(988);
     data_out(4843) <= data_in(990);
     data_out(4844) <= data_in(992);
     data_out(4845) <= data_in(995);
     data_out(4846) <= data_in(998);
     data_out(4847) <= data_in(1000);
     data_out(4848) <= data_in(1003);
     data_out(4849) <= data_in(1006);
     data_out(4850) <= data_in(1011);
     data_out(4851) <= data_in(1012);
     data_out(4852) <= data_in(1020);
     data_out(4853) <= data_in(1022);
     data_out(4854) <= data_in(1026);
     data_out(4855) <= data_in(1030);
     data_out(4856) <= data_in(1034);
     data_out(4857) <= data_in(1035);
     data_out(4858) <= data_in(1039);
     data_out(4859) <= data_in(1044);
     data_out(4860) <= data_in(1046);
     data_out(4861) <= data_in(1049);
     data_out(4862) <= data_in(1069);
     data_out(4863) <= data_in(1072);
     data_out(4864) <= data_in(1073);
     data_out(4865) <= data_in(1076);
     data_out(4866) <= data_in(1077);
     data_out(4867) <= data_in(1082);
     data_out(4868) <= data_in(1090);
     data_out(4869) <= data_in(1091);
     data_out(4870) <= data_in(1092);
     data_out(4871) <= data_in(1097);
     data_out(4872) <= data_in(1098);
     data_out(4873) <= data_in(1101);
     data_out(4874) <= data_in(1104);
     data_out(4875) <= data_in(1106);
     data_out(4876) <= data_in(1115);
     data_out(4877) <= data_in(1117);
     data_out(4878) <= data_in(1118);
     data_out(4879) <= data_in(1124);
     data_out(4880) <= data_in(1125);
     data_out(4881) <= data_in(1127);
     data_out(4882) <= data_in(1129);
     data_out(4883) <= data_in(1130);
     data_out(4884) <= data_in(1131);
     data_out(4885) <= data_in(1134);
     data_out(4886) <= data_in(1135);
     data_out(4887) <= data_in(1136);
     data_out(4888) <= data_in(1137);
     data_out(4889) <= data_in(1138);
     data_out(4890) <= data_in(1139);
     data_out(4891) <= data_in(1142);
     data_out(4892) <= data_in(1144);
     data_out(4893) <= data_in(1146);
     data_out(4894) <= data_in(1147);
     data_out(4895) <= data_in(1150);
     data_out(4896) <= data_in(1151);
     data_out(4897) <= data_in(1153);
     data_out(4898) <= data_in(1154);
     data_out(4899) <= data_in(1155);
     data_out(4900) <= data_in(1156);
     data_out(4901) <= data_in(1157);
     data_out(4902) <= data_in(1160);
     data_out(4903) <= data_in(1165);
     data_out(4904) <= data_in(1166);
     data_out(4905) <= data_in(1167);
     data_out(4906) <= data_in(1170);
     data_out(4907) <= data_in(1175);
     data_out(4908) <= data_in(1179);
     data_out(4909) <= data_in(1182);
     data_out(4910) <= data_in(1184);
     data_out(4911) <= data_in(1186);
     data_out(4912) <= data_in(1194);
     data_out(4913) <= data_in(1200);
     data_out(4914) <= data_in(1201);
     data_out(4915) <= data_in(1202);
     data_out(4916) <= data_in(1204);
     data_out(4917) <= data_in(1206);
     data_out(4918) <= data_in(1209);
     data_out(4919) <= data_in(1214);
     data_out(4920) <= data_in(1221);
     data_out(4921) <= data_in(1222);
     data_out(4922) <= data_in(1231);
     data_out(4923) <= data_in(1234);
     data_out(4924) <= data_in(1235);
     data_out(4925) <= data_in(1236);
     data_out(4926) <= data_in(1238);
     data_out(4927) <= data_in(1243);
     data_out(4928) <= data_in(1245);
     data_out(4929) <= data_in(1246);
     data_out(4930) <= data_in(1248);
     data_out(4931) <= data_in(1253);
     data_out(4932) <= data_in(1259);
     data_out(4933) <= data_in(1264);
     data_out(4934) <= data_in(1265);
     data_out(4935) <= data_in(1266);
     data_out(4936) <= data_in(1268);
     data_out(4937) <= data_in(1270);
     data_out(4938) <= data_in(1272);
     data_out(4939) <= data_in(1275);
     data_out(4940) <= data_in(1276);
     data_out(4941) <= data_in(1278);
     data_out(4942) <= data_in(1282);
     data_out(4943) <= data_in(1284);
     data_out(4944) <= data_in(1288);
     data_out(4945) <= data_in(1289);
     data_out(4946) <= data_in(1290);
     data_out(4947) <= data_in(1292);
     data_out(4948) <= data_in(1299);
     data_out(4949) <= data_in(1300);
     data_out(4950) <= data_in(1301);
     data_out(4951) <= data_in(1303);
     data_out(4952) <= data_in(1306);
     data_out(4953) <= data_in(1312);
     data_out(4954) <= data_in(1315);
     data_out(4955) <= data_in(1318);
     data_out(4956) <= data_in(1319);
     data_out(4957) <= data_in(1321);
     data_out(4958) <= data_in(1322);
     data_out(4959) <= data_in(1324);
     data_out(4960) <= data_in(1325);
     data_out(4961) <= data_in(1334);
     data_out(4962) <= data_in(1335);
     data_out(4963) <= data_in(1336);
     data_out(4964) <= data_in(1340);
     data_out(4965) <= data_in(1342);
     data_out(4966) <= data_in(1346);
     data_out(4967) <= data_in(1348);
     data_out(4968) <= data_in(1351);
     data_out(4969) <= data_in(1353);
     data_out(4970) <= data_in(1355);
     data_out(4971) <= data_in(1356);
     data_out(4972) <= data_in(1357);
     data_out(4973) <= data_in(1367);
     data_out(4974) <= data_in(1368);
     data_out(4975) <= data_in(1371);
     data_out(4976) <= data_in(1373);
     data_out(4977) <= data_in(1376);
     data_out(4978) <= data_in(1377);
     data_out(4979) <= data_in(1380);
     data_out(4980) <= data_in(1383);
     data_out(4981) <= data_in(1387);
     data_out(4982) <= data_in(1388);
     data_out(4983) <= data_in(1391);
     data_out(4984) <= data_in(1393);
     data_out(4985) <= data_in(1394);
     data_out(4986) <= data_in(1396);
     data_out(4987) <= data_in(1397);
     data_out(4988) <= data_in(1398);
     data_out(4989) <= data_in(1400);
     data_out(4990) <= data_in(1404);
     data_out(4991) <= data_in(1405);
     data_out(4992) <= data_in(1410);
     data_out(4993) <= data_in(1411);
     data_out(4994) <= data_in(1413);
     data_out(4995) <= data_in(1417);
     data_out(4996) <= data_in(1420);
     data_out(4997) <= data_in(1421);
     data_out(4998) <= data_in(1427);
     data_out(4999) <= data_in(1433);
     data_out(5000) <= data_in(1434);
     data_out(5001) <= data_in(1435);
     data_out(5002) <= data_in(1437);
     data_out(5003) <= data_in(1442);
     data_out(5004) <= data_in(1443);
     data_out(5005) <= data_in(1448);
     data_out(5006) <= data_in(1449);
     data_out(5007) <= data_in(1452);
     data_out(5008) <= data_in(1454);
     data_out(5009) <= data_in(1456);
     data_out(5010) <= data_in(1463);
     data_out(5011) <= data_in(1464);
     data_out(5012) <= data_in(1467);
     data_out(5013) <= data_in(1471);
     data_out(5014) <= data_in(1472);
     data_out(5015) <= data_in(1473);
     data_out(5016) <= data_in(1477);
     data_out(5017) <= data_in(1479);
     data_out(5018) <= data_in(1484);
     data_out(5019) <= data_in(1493);
     data_out(5020) <= data_in(1495);
     data_out(5021) <= data_in(1498);
     data_out(5022) <= data_in(1500);
     data_out(5023) <= data_in(1502);
     data_out(5024) <= data_in(1503);
     data_out(5025) <= data_in(1519);
     data_out(5026) <= data_in(1520);
     data_out(5027) <= data_in(1523);
     data_out(5028) <= data_in(1525);
     data_out(5029) <= data_in(1527);
     data_out(5030) <= data_in(1528);
     data_out(5031) <= data_in(1531);
     data_out(5032) <= data_in(1539);
     data_out(5033) <= data_in(1540);
     data_out(5034) <= data_in(1547);
     data_out(5035) <= data_in(1549);
     data_out(5036) <= data_in(1552);
     data_out(5037) <= data_in(1556);
     data_out(5038) <= data_in(1563);
     data_out(5039) <= data_in(1564);
     data_out(5040) <= data_in(1566);
     data_out(5041) <= data_in(1568);
     data_out(5042) <= data_in(1570);
     data_out(5043) <= data_in(1573);
     data_out(5044) <= data_in(1576);
     data_out(5045) <= data_in(1581);
     data_out(5046) <= data_in(1582);
     data_out(5047) <= data_in(1583);
     data_out(5048) <= data_in(1585);
     data_out(5049) <= data_in(1591);
     data_out(5050) <= data_in(1595);
     data_out(5051) <= data_in(1602);
     data_out(5052) <= data_in(1605);
     data_out(5053) <= data_in(1609);
     data_out(5054) <= data_in(1612);
     data_out(5055) <= data_in(1617);
     data_out(5056) <= data_in(1618);
     data_out(5057) <= data_in(1619);
     data_out(5058) <= data_in(1621);
     data_out(5059) <= data_in(1623);
     data_out(5060) <= data_in(1627);
     data_out(5061) <= data_in(1630);
     data_out(5062) <= data_in(1631);
     data_out(5063) <= data_in(1632);
     data_out(5064) <= data_in(1633);
     data_out(5065) <= data_in(1635);
     data_out(5066) <= data_in(1642);
     data_out(5067) <= data_in(1644);
     data_out(5068) <= data_in(1648);
     data_out(5069) <= data_in(1650);
     data_out(5070) <= data_in(1652);
     data_out(5071) <= data_in(1653);
     data_out(5072) <= data_in(1654);
     data_out(5073) <= data_in(1656);
     data_out(5074) <= data_in(1657);
     data_out(5075) <= data_in(1661);
     data_out(5076) <= data_in(1662);
     data_out(5077) <= data_in(1663);
     data_out(5078) <= data_in(1665);
     data_out(5079) <= data_in(1669);
     data_out(5080) <= data_in(1672);
     data_out(5081) <= data_in(1673);
     data_out(5082) <= data_in(1677);
     data_out(5083) <= data_in(1679);
     data_out(5084) <= data_in(1680);
     data_out(5085) <= data_in(1683);
     data_out(5086) <= data_in(1690);
     data_out(5087) <= data_in(1692);
     data_out(5088) <= data_in(1693);
     data_out(5089) <= data_in(1696);
     data_out(5090) <= data_in(1698);
     data_out(5091) <= data_in(1702);
     data_out(5092) <= data_in(1704);
     data_out(5093) <= data_in(1706);
     data_out(5094) <= data_in(1707);
     data_out(5095) <= data_in(1708);
     data_out(5096) <= data_in(1709);
     data_out(5097) <= data_in(1715);
     data_out(5098) <= data_in(1716);
     data_out(5099) <= data_in(1718);
     data_out(5100) <= data_in(1722);
     data_out(5101) <= data_in(1724);
     data_out(5102) <= data_in(1732);
     data_out(5103) <= data_in(1733);
     data_out(5104) <= data_in(1735);
     data_out(5105) <= data_in(1736);
     data_out(5106) <= data_in(1738);
     data_out(5107) <= data_in(1739);
     data_out(5108) <= data_in(1745);
     data_out(5109) <= data_in(1746);
     data_out(5110) <= data_in(1749);
     data_out(5111) <= data_in(1751);
     data_out(5112) <= data_in(1752);
     data_out(5113) <= data_in(1753);
     data_out(5114) <= data_in(1755);
     data_out(5115) <= data_in(1756);
     data_out(5116) <= data_in(1758);
     data_out(5117) <= data_in(1759);
     data_out(5118) <= data_in(1760);
     data_out(5119) <= data_in(1761);
     data_out(5120) <= data_in(1765);
     data_out(5121) <= data_in(1769);
     data_out(5122) <= data_in(1771);
     data_out(5123) <= data_in(1775);
     data_out(5124) <= data_in(1776);
     data_out(5125) <= data_in(1778);
     data_out(5126) <= data_in(1785);
     data_out(5127) <= data_in(1787);
     data_out(5128) <= data_in(1791);
     data_out(5129) <= data_in(1792);
     data_out(5130) <= data_in(1798);
     data_out(5131) <= data_in(1799);
     data_out(5132) <= data_in(1801);
     data_out(5133) <= data_in(1802);
     data_out(5134) <= data_in(1808);
     data_out(5135) <= data_in(1814);
     data_out(5136) <= data_in(1816);
     data_out(5137) <= data_in(1819);
     data_out(5138) <= data_in(1822);
     data_out(5139) <= data_in(1823);
     data_out(5140) <= data_in(1830);
     data_out(5141) <= data_in(1831);
     data_out(5142) <= data_in(1832);
     data_out(5143) <= data_in(1834);
     data_out(5144) <= data_in(1838);
     data_out(5145) <= data_in(1840);
     data_out(5146) <= data_in(1845);
     data_out(5147) <= data_in(1846);
     data_out(5148) <= data_in(1849);
     data_out(5149) <= data_in(1851);
     data_out(5150) <= data_in(1856);
     data_out(5151) <= data_in(1857);
     data_out(5152) <= data_in(1861);
     data_out(5153) <= data_in(1863);
     data_out(5154) <= data_in(1865);
     data_out(5155) <= data_in(1866);
     data_out(5156) <= data_in(1868);
     data_out(5157) <= data_in(1870);
     data_out(5158) <= data_in(1871);
     data_out(5159) <= data_in(1874);
     data_out(5160) <= data_in(1880);
     data_out(5161) <= data_in(1881);
     data_out(5162) <= data_in(1882);
     data_out(5163) <= data_in(1888);
     data_out(5164) <= data_in(1894);
     data_out(5165) <= data_in(1901);
     data_out(5166) <= data_in(1903);
     data_out(5167) <= data_in(1905);
     data_out(5168) <= data_in(1909);
     data_out(5169) <= data_in(1920);
     data_out(5170) <= data_in(1923);
     data_out(5171) <= data_in(1927);
     data_out(5172) <= data_in(1929);
     data_out(5173) <= data_in(1932);
     data_out(5174) <= data_in(1940);
     data_out(5175) <= data_in(1942);
     data_out(5176) <= data_in(1943);
     data_out(5177) <= data_in(1944);
     data_out(5178) <= data_in(1946);
     data_out(5179) <= data_in(1949);
     data_out(5180) <= data_in(1953);
     data_out(5181) <= data_in(1954);
     data_out(5182) <= data_in(1956);
     data_out(5183) <= data_in(1962);
     data_out(5184) <= data_in(1963);
     data_out(5185) <= data_in(1969);
     data_out(5186) <= data_in(1972);
     data_out(5187) <= data_in(1973);
     data_out(5188) <= data_in(1978);
     data_out(5189) <= data_in(1983);
     data_out(5190) <= data_in(1988);
     data_out(5191) <= data_in(1991);
     data_out(5192) <= data_in(1997);
     data_out(5193) <= data_in(1998);
     data_out(5194) <= data_in(2002);
     data_out(5195) <= data_in(2003);
     data_out(5196) <= data_in(2009);
     data_out(5197) <= data_in(2013);
     data_out(5198) <= data_in(2014);
     data_out(5199) <= data_in(2015);
     data_out(5200) <= data_in(2016);
     data_out(5201) <= data_in(2017);
     data_out(5202) <= data_in(2019);
     data_out(5203) <= data_in(2023);
     data_out(5204) <= data_in(2025);
     data_out(5205) <= data_in(2027);
     data_out(5206) <= data_in(2029);
     data_out(5207) <= data_in(2030);
     data_out(5208) <= data_in(2031);
     data_out(5209) <= data_in(2032);
     data_out(5210) <= data_in(2033);
     data_out(5211) <= data_in(2043);
     data_out(5212) <= data_in(2045);
     data_out(5213) <= data_in(2047);
     data_out(5214) <= data_in(2048);
     data_out(5215) <= data_in(2050);
     data_out(5216) <= data_in(2052);
     data_out(5217) <= data_in(2054);
     data_out(5218) <= data_in(2055);
     data_out(5219) <= data_in(2056);
     data_out(5220) <= data_in(2061);
     data_out(5221) <= data_in(2063);
     data_out(5222) <= data_in(2065);
     data_out(5223) <= data_in(2067);
     data_out(5224) <= data_in(2068);
     data_out(5225) <= data_in(2070);
     data_out(5226) <= data_in(2074);
     data_out(5227) <= data_in(2078);
     data_out(5228) <= data_in(2083);
     data_out(5229) <= data_in(2084);
     data_out(5230) <= data_in(2090);
     data_out(5231) <= data_in(2092);
     data_out(5232) <= data_in(2094);
     data_out(5233) <= data_in(2095);
     data_out(5234) <= data_in(2104);
     data_out(5235) <= data_in(2109);
     data_out(5236) <= data_in(2110);
     data_out(5237) <= data_in(2112);
     data_out(5238) <= data_in(2113);
     data_out(5239) <= data_in(2116);
     data_out(5240) <= data_in(2117);
     data_out(5241) <= data_in(2120);
     data_out(5242) <= data_in(2122);
     data_out(5243) <= data_in(2126);
     data_out(5244) <= data_in(2127);
     data_out(5245) <= data_in(2130);
     data_out(5246) <= data_in(2132);
     data_out(5247) <= data_in(2137);
     data_out(5248) <= data_in(2144);
     data_out(5249) <= data_in(2147);
     data_out(5250) <= data_in(2151);
     data_out(5251) <= data_in(2155);
     data_out(5252) <= data_in(2156);
     data_out(5253) <= data_in(2157);
     data_out(5254) <= data_in(2159);
     data_out(5255) <= data_in(2160);
     data_out(5256) <= data_in(2161);
     data_out(5257) <= data_in(2162);
     data_out(5258) <= data_in(2166);
     data_out(5259) <= data_in(2168);
     data_out(5260) <= data_in(2169);
     data_out(5261) <= data_in(2171);
     data_out(5262) <= data_in(2181);
     data_out(5263) <= data_in(2182);
     data_out(5264) <= data_in(2188);
     data_out(5265) <= data_in(2190);
     data_out(5266) <= data_in(2192);
     data_out(5267) <= data_in(2196);
     data_out(5268) <= data_in(2198);
     data_out(5269) <= data_in(2199);
     data_out(5270) <= data_in(2201);
     data_out(5271) <= data_in(2202);
     data_out(5272) <= data_in(2203);
     data_out(5273) <= data_in(2205);
     data_out(5274) <= data_in(2206);
     data_out(5275) <= data_in(2207);
     data_out(5276) <= data_in(2208);
     data_out(5277) <= data_in(2209);
     data_out(5278) <= data_in(2210);
     data_out(5279) <= data_in(2215);
     data_out(5280) <= data_in(2216);
     data_out(5281) <= data_in(2219);
     data_out(5282) <= data_in(2220);
     data_out(5283) <= data_in(2222);
     data_out(5284) <= data_in(2229);
     data_out(5285) <= data_in(2233);
     data_out(5286) <= data_in(2239);
     data_out(5287) <= data_in(2240);
     data_out(5288) <= data_in(2246);
     data_out(5289) <= data_in(2249);
     data_out(5290) <= data_in(2250);
     data_out(5291) <= data_in(2251);
     data_out(5292) <= data_in(2257);
     data_out(5293) <= data_in(2258);
     data_out(5294) <= data_in(2260);
     data_out(5295) <= data_in(2261);
     data_out(5296) <= data_in(2263);
     data_out(5297) <= data_in(2269);
     data_out(5298) <= data_in(2271);
     data_out(5299) <= data_in(2276);
     data_out(5300) <= data_in(2282);
     data_out(5301) <= data_in(2286);
     data_out(5302) <= data_in(2288);
     data_out(5303) <= data_in(2292);
     data_out(5304) <= data_in(2295);
     data_out(5305) <= data_in(2298);
     data_out(5306) <= data_in(2300);
     data_out(5307) <= data_in(2301);
     data_out(5308) <= data_in(2302);
     data_out(5309) <= data_in(2303);
     data_out(5310) <= data_in(2310);
     data_out(5311) <= data_in(2311);
     data_out(5312) <= data_in(2316);
     data_out(5313) <= data_in(2317);
     data_out(5314) <= data_in(2319);
     data_out(5315) <= data_in(2321);
     data_out(5316) <= data_in(2325);
     data_out(5317) <= data_in(2327);
     data_out(5318) <= data_in(2330);
     data_out(5319) <= data_in(2335);
     data_out(5320) <= data_in(2340);
     data_out(5321) <= data_in(2342);
     data_out(5322) <= data_in(2343);
     data_out(5323) <= data_in(2349);
     data_out(5324) <= data_in(2350);
     data_out(5325) <= data_in(2354);
     data_out(5326) <= data_in(2356);
     data_out(5327) <= data_in(2357);
     data_out(5328) <= data_in(2360);
     data_out(5329) <= data_in(2363);
     data_out(5330) <= data_in(2364);
     data_out(5331) <= data_in(2367);
     data_out(5332) <= data_in(2369);
     data_out(5333) <= data_in(2374);
     data_out(5334) <= data_in(2380);
     data_out(5335) <= data_in(2382);
     data_out(5336) <= data_in(2383);
     data_out(5337) <= data_in(2384);
     data_out(5338) <= data_in(2387);
     data_out(5339) <= data_in(2388);
     data_out(5340) <= data_in(2392);
     data_out(5341) <= data_in(2393);
     data_out(5342) <= data_in(2398);
     data_out(5343) <= data_in(2400);
     data_out(5344) <= data_in(2401);
     data_out(5345) <= data_in(2402);
     data_out(5346) <= data_in(2403);
     data_out(5347) <= data_in(2405);
     data_out(5348) <= data_in(2412);
     data_out(5349) <= data_in(2413);
     data_out(5350) <= data_in(2415);
     data_out(5351) <= data_in(2419);
     data_out(5352) <= data_in(2420);
     data_out(5353) <= data_in(2422);
     data_out(5354) <= data_in(2424);
     data_out(5355) <= data_in(2426);
     data_out(5356) <= data_in(2431);
     data_out(5357) <= data_in(2432);
     data_out(5358) <= data_in(2436);
     data_out(5359) <= data_in(2439);
     data_out(5360) <= data_in(2443);
     data_out(5361) <= data_in(2446);
     data_out(5362) <= data_in(2447);
     data_out(5363) <= data_in(2451);
     data_out(5364) <= data_in(2453);
     data_out(5365) <= data_in(2456);
     data_out(5366) <= data_in(2461);
     data_out(5367) <= data_in(2462);
     data_out(5368) <= data_in(2464);
     data_out(5369) <= data_in(2465);
     data_out(5370) <= data_in(2466);
     data_out(5371) <= data_in(2470);
     data_out(5372) <= data_in(2472);
     data_out(5373) <= data_in(2474);
     data_out(5374) <= data_in(2475);
     data_out(5375) <= data_in(2477);
     data_out(5376) <= data_in(2479);
     data_out(5377) <= data_in(2481);
     data_out(5378) <= data_in(2482);
     data_out(5379) <= data_in(2484);
     data_out(5380) <= data_in(2487);
     data_out(5381) <= data_in(2488);
     data_out(5382) <= data_in(2492);
     data_out(5383) <= data_in(2493);
     data_out(5384) <= data_in(2494);
     data_out(5385) <= data_in(2495);
     data_out(5386) <= data_in(2498);
     data_out(5387) <= data_in(2505);
     data_out(5388) <= data_in(2506);
     data_out(5389) <= data_in(2509);
     data_out(5390) <= data_in(2510);
     data_out(5391) <= data_in(2511);
     data_out(5392) <= data_in(2512);
     data_out(5393) <= data_in(2517);
     data_out(5394) <= data_in(2519);
     data_out(5395) <= data_in(2525);
     data_out(5396) <= data_in(2526);
     data_out(5397) <= data_in(2527);
     data_out(5398) <= data_in(2531);
     data_out(5399) <= data_in(2535);
     data_out(5400) <= data_in(2539);
     data_out(5401) <= data_in(2540);
     data_out(5402) <= data_in(2543);
     data_out(5403) <= data_in(2551);
     data_out(5404) <= data_in(2552);
     data_out(5405) <= data_in(2556);
     data_out(5406) <= data_in(2558);
     data_out(5407) <= data_in(2560);
     data_out(5408) <= data_in(2563);
     data_out(5409) <= data_in(2564);
     data_out(5410) <= data_in(2566);
     data_out(5411) <= data_in(2568);
     data_out(5412) <= data_in(2569);
     data_out(5413) <= data_in(2571);
     data_out(5414) <= data_in(2572);
     data_out(5415) <= data_in(2577);
     data_out(5416) <= data_in(2578);
     data_out(5417) <= data_in(2590);
     data_out(5418) <= data_in(2591);
     data_out(5419) <= data_in(2597);
     data_out(5420) <= data_in(2599);
     data_out(5421) <= data_in(2600);
     data_out(5422) <= data_in(2602);
     data_out(5423) <= data_in(2603);
     data_out(5424) <= data_in(2604);
     data_out(5425) <= data_in(2605);
     data_out(5426) <= data_in(2606);
     data_out(5427) <= data_in(2609);
     data_out(5428) <= data_in(2613);
     data_out(5429) <= data_in(2616);
     data_out(5430) <= data_in(2620);
     data_out(5431) <= data_in(2627);
     data_out(5432) <= data_in(2630);
     data_out(5433) <= data_in(2631);
     data_out(5434) <= data_in(2636);
     data_out(5435) <= data_in(2637);
     data_out(5436) <= data_in(2639);
     data_out(5437) <= data_in(2641);
     data_out(5438) <= data_in(2648);
     data_out(5439) <= data_in(2649);
     data_out(5440) <= data_in(2650);
     data_out(5441) <= data_in(2658);
     data_out(5442) <= data_in(2659);
     data_out(5443) <= data_in(2665);
     data_out(5444) <= data_in(2675);
     data_out(5445) <= data_in(2680);
     data_out(5446) <= data_in(2681);
     data_out(5447) <= data_in(2685);
     data_out(5448) <= data_in(2687);
     data_out(5449) <= data_in(2688);
     data_out(5450) <= data_in(2694);
     data_out(5451) <= data_in(2695);
     data_out(5452) <= data_in(2704);
     data_out(5453) <= data_in(2706);
     data_out(5454) <= data_in(2708);
     data_out(5455) <= data_in(2709);
     data_out(5456) <= data_in(2718);
     data_out(5457) <= data_in(2719);
     data_out(5458) <= data_in(2720);
     data_out(5459) <= data_in(2727);
     data_out(5460) <= data_in(2728);
     data_out(5461) <= data_in(2729);
     data_out(5462) <= data_in(2734);
     data_out(5463) <= data_in(2735);
     data_out(5464) <= data_in(2736);
     data_out(5465) <= data_in(2737);
     data_out(5466) <= data_in(2740);
     data_out(5467) <= data_in(2744);
     data_out(5468) <= data_in(2745);
     data_out(5469) <= data_in(2747);
     data_out(5470) <= data_in(2754);
     data_out(5471) <= data_in(2756);
     data_out(5472) <= data_in(2757);
     data_out(5473) <= data_in(2758);
     data_out(5474) <= data_in(2763);
     data_out(5475) <= data_in(2766);
     data_out(5476) <= data_in(2768);
     data_out(5477) <= data_in(2769);
     data_out(5478) <= data_in(2772);
     data_out(5479) <= data_in(2775);
     data_out(5480) <= data_in(2777);
     data_out(5481) <= data_in(2781);
     data_out(5482) <= data_in(2788);
     data_out(5483) <= data_in(2790);
     data_out(5484) <= data_in(2793);
     data_out(5485) <= data_in(2794);
     data_out(5486) <= data_in(2795);
     data_out(5487) <= data_in(2797);
     data_out(5488) <= data_in(2798);
     data_out(5489) <= data_in(2799);
     data_out(5490) <= data_in(2800);
     data_out(5491) <= data_in(2802);
     data_out(5492) <= data_in(2806);
     data_out(5493) <= data_in(2807);
     data_out(5494) <= data_in(2813);
     data_out(5495) <= data_in(2815);
     data_out(5496) <= data_in(2817);
     data_out(5497) <= data_in(2818);
     data_out(5498) <= data_in(2819);
     data_out(5499) <= data_in(2820);
     data_out(5500) <= data_in(2825);
     data_out(5501) <= data_in(2827);
     data_out(5502) <= data_in(2828);
     data_out(5503) <= data_in(2834);
     data_out(5504) <= data_in(2835);
     data_out(5505) <= data_in(2836);
     data_out(5506) <= data_in(2838);
     data_out(5507) <= data_in(2840);
     data_out(5508) <= data_in(2845);
     data_out(5509) <= data_in(2846);
     data_out(5510) <= data_in(2847);
     data_out(5511) <= data_in(2851);
     data_out(5512) <= data_in(2858);
     data_out(5513) <= data_in(2859);
     data_out(5514) <= data_in(2861);
     data_out(5515) <= data_in(2866);
     data_out(5516) <= data_in(2868);
     data_out(5517) <= data_in(2869);
     data_out(5518) <= data_in(2870);
     data_out(5519) <= data_in(2871);
     data_out(5520) <= data_in(2872);
     data_out(5521) <= data_in(2877);
     data_out(5522) <= data_in(2882);
     data_out(5523) <= data_in(2883);
     data_out(5524) <= data_in(2886);
     data_out(5525) <= data_in(2891);
     data_out(5526) <= data_in(2893);
     data_out(5527) <= data_in(2898);
     data_out(5528) <= data_in(2902);
     data_out(5529) <= data_in(2903);
     data_out(5530) <= data_in(2904);
     data_out(5531) <= data_in(2905);
     data_out(5532) <= data_in(2906);
     data_out(5533) <= data_in(2909);
     data_out(5534) <= data_in(2911);
     data_out(5535) <= data_in(2914);
     data_out(5536) <= data_in(2920);
     data_out(5537) <= data_in(2922);
     data_out(5538) <= data_in(2928);
     data_out(5539) <= data_in(2935);
     data_out(5540) <= data_in(2938);
     data_out(5541) <= data_in(2942);
     data_out(5542) <= data_in(2943);
     data_out(5543) <= data_in(2946);
     data_out(5544) <= data_in(2951);
     data_out(5545) <= data_in(2952);
     data_out(5546) <= data_in(2955);
     data_out(5547) <= data_in(2958);
     data_out(5548) <= data_in(2966);
     data_out(5549) <= data_in(2969);
     data_out(5550) <= data_in(2971);
     data_out(5551) <= data_in(2978);
     data_out(5552) <= data_in(2979);
     data_out(5553) <= data_in(2980);
     data_out(5554) <= data_in(2982);
     data_out(5555) <= data_in(2984);
     data_out(5556) <= data_in(2986);
     data_out(5557) <= data_in(2992);
     data_out(5558) <= data_in(2996);
     data_out(5559) <= data_in(3000);
     data_out(5560) <= data_in(3001);
     data_out(5561) <= data_in(3002);
     data_out(5562) <= data_in(3008);
     data_out(5563) <= data_in(3009);
     data_out(5564) <= data_in(3010);
     data_out(5565) <= data_in(3013);
     data_out(5566) <= data_in(3014);
     data_out(5567) <= data_in(3017);
     data_out(5568) <= data_in(3019);
     data_out(5569) <= data_in(3023);
     data_out(5570) <= data_in(3024);
     data_out(5571) <= data_in(3028);
     data_out(5572) <= data_in(3036);
     data_out(5573) <= data_in(3040);
     data_out(5574) <= data_in(3043);
     data_out(5575) <= data_in(3045);
     data_out(5576) <= data_in(3047);
     data_out(5577) <= data_in(3048);
     data_out(5578) <= data_in(3051);
     data_out(5579) <= data_in(3052);
     data_out(5580) <= data_in(3056);
     data_out(5581) <= data_in(3058);
     data_out(5582) <= data_in(3062);
     data_out(5583) <= data_in(3067);
     data_out(5584) <= data_in(3068);
     data_out(5585) <= data_in(3069);
     data_out(5586) <= data_in(3070);
     data_out(5587) <= data_in(3074);
     data_out(5588) <= data_in(3076);
     data_out(5589) <= data_in(3078);
     data_out(5590) <= data_in(3079);
     data_out(5591) <= data_in(3082);
     data_out(5592) <= data_in(3087);
     data_out(5593) <= data_in(3089);
     data_out(5594) <= data_in(3096);
     data_out(5595) <= data_in(3098);
     data_out(5596) <= data_in(3099);
     data_out(5597) <= data_in(3102);
     data_out(5598) <= data_in(3105);
     data_out(5599) <= data_in(3110);
     data_out(5600) <= data_in(3111);
     data_out(5601) <= data_in(3112);
     data_out(5602) <= data_in(3113);
     data_out(5603) <= data_in(3114);
     data_out(5604) <= data_in(3117);
     data_out(5605) <= data_in(3118);
     data_out(5606) <= data_in(3120);
     data_out(5607) <= data_in(3121);
     data_out(5608) <= data_in(3122);
     data_out(5609) <= data_in(3125);
     data_out(5610) <= data_in(3130);
     data_out(5611) <= data_in(3131);
     data_out(5612) <= data_in(3132);
     data_out(5613) <= data_in(3134);
     data_out(5614) <= data_in(3137);
     data_out(5615) <= data_in(3142);
     data_out(5616) <= data_in(3144);
     data_out(5617) <= data_in(3148);
     data_out(5618) <= data_in(3152);
     data_out(5619) <= data_in(3155);
     data_out(5620) <= data_in(3156);
     data_out(5621) <= data_in(3158);
     data_out(5622) <= data_in(3159);
     data_out(5623) <= data_in(3161);
     data_out(5624) <= data_in(3163);
     data_out(5625) <= data_in(3168);
     data_out(5626) <= data_in(3171);
     data_out(5627) <= data_in(3173);
     data_out(5628) <= data_in(3178);
     data_out(5629) <= data_in(3185);
     data_out(5630) <= data_in(3186);
     data_out(5631) <= data_in(3187);
     data_out(5632) <= data_in(3190);
     data_out(5633) <= data_in(3192);
     data_out(5634) <= data_in(3193);
     data_out(5635) <= data_in(3195);
     data_out(5636) <= data_in(3200);
     data_out(5637) <= data_in(3201);
     data_out(5638) <= data_in(3207);
     data_out(5639) <= data_in(3211);
     data_out(5640) <= data_in(3216);
     data_out(5641) <= data_in(3219);
     data_out(5642) <= data_in(3221);
     data_out(5643) <= data_in(3224);
     data_out(5644) <= data_in(3225);
     data_out(5645) <= data_in(3230);
     data_out(5646) <= data_in(3231);
     data_out(5647) <= data_in(3233);
     data_out(5648) <= data_in(3237);
     data_out(5649) <= data_in(3238);
     data_out(5650) <= data_in(3239);
     data_out(5651) <= data_in(3241);
     data_out(5652) <= data_in(3243);
     data_out(5653) <= data_in(3244);
     data_out(5654) <= data_in(3248);
     data_out(5655) <= data_in(3250);
     data_out(5656) <= data_in(3253);
     data_out(5657) <= data_in(3256);
     data_out(5658) <= data_in(3257);
     data_out(5659) <= data_in(3261);
     data_out(5660) <= data_in(3262);
     data_out(5661) <= data_in(3265);
     data_out(5662) <= data_in(3269);
     data_out(5663) <= data_in(3272);
     data_out(5664) <= data_in(3273);
     data_out(5665) <= data_in(3276);
     data_out(5666) <= data_in(3280);
     data_out(5667) <= data_in(3281);
     data_out(5668) <= data_in(3283);
     data_out(5669) <= data_in(3284);
     data_out(5670) <= data_in(3288);
     data_out(5671) <= data_in(3289);
     data_out(5672) <= data_in(3290);
     data_out(5673) <= data_in(3291);
     data_out(5674) <= data_in(3294);
     data_out(5675) <= data_in(3299);
     data_out(5676) <= data_in(3311);
     data_out(5677) <= data_in(3317);
     data_out(5678) <= data_in(3320);
     data_out(5679) <= data_in(3326);
     data_out(5680) <= data_in(3336);
     data_out(5681) <= data_in(3337);
     data_out(5682) <= data_in(3341);
     data_out(5683) <= data_in(3344);
     data_out(5684) <= data_in(3346);
     data_out(5685) <= data_in(3348);
     data_out(5686) <= data_in(3350);
     data_out(5687) <= data_in(3351);
     data_out(5688) <= data_in(3352);
     data_out(5689) <= data_in(3354);
     data_out(5690) <= data_in(3355);
     data_out(5691) <= data_in(3357);
     data_out(5692) <= data_in(3362);
     data_out(5693) <= data_in(3366);
     data_out(5694) <= data_in(3367);
     data_out(5695) <= data_in(3368);
     data_out(5696) <= data_in(3370);
     data_out(5697) <= data_in(3371);
     data_out(5698) <= data_in(3376);
     data_out(5699) <= data_in(3378);
     data_out(5700) <= data_in(3380);
     data_out(5701) <= data_in(3381);
     data_out(5702) <= data_in(3382);
     data_out(5703) <= data_in(3385);
     data_out(5704) <= data_in(3388);
     data_out(5705) <= data_in(3392);
     data_out(5706) <= data_in(3396);
     data_out(5707) <= data_in(3399);
     data_out(5708) <= data_in(3401);
     data_out(5709) <= data_in(3407);
     data_out(5710) <= data_in(3408);
     data_out(5711) <= data_in(3418);
     data_out(5712) <= data_in(3420);
     data_out(5713) <= data_in(3423);
     data_out(5714) <= data_in(3430);
     data_out(5715) <= data_in(3431);
     data_out(5716) <= data_in(3432);
     data_out(5717) <= data_in(3434);
     data_out(5718) <= data_in(3439);
     data_out(5719) <= data_in(3443);
     data_out(5720) <= data_in(3444);
     data_out(5721) <= data_in(3445);
     data_out(5722) <= data_in(3446);
     data_out(5723) <= data_in(3447);
     data_out(5724) <= data_in(3449);
     data_out(5725) <= data_in(3451);
     data_out(5726) <= data_in(3452);
     data_out(5727) <= data_in(3453);
     data_out(5728) <= data_in(3454);
     data_out(5729) <= data_in(3457);
     data_out(5730) <= data_in(3458);
     data_out(5731) <= data_in(3460);
     data_out(5732) <= data_in(3461);
     data_out(5733) <= data_in(3465);
     data_out(5734) <= data_in(3467);
     data_out(5735) <= data_in(3469);
     data_out(5736) <= data_in(3471);
     data_out(5737) <= data_in(3473);
     data_out(5738) <= data_in(3476);
     data_out(5739) <= data_in(3480);
     data_out(5740) <= data_in(3481);
     data_out(5741) <= data_in(3482);
     data_out(5742) <= data_in(3483);
     data_out(5743) <= data_in(3487);
     data_out(5744) <= data_in(3489);
     data_out(5745) <= data_in(3490);
     data_out(5746) <= data_in(3493);
     data_out(5747) <= data_in(3496);
     data_out(5748) <= data_in(3499);
     data_out(5749) <= data_in(3500);
     data_out(5750) <= data_in(3501);
     data_out(5751) <= data_in(3502);
     data_out(5752) <= data_in(3505);
     data_out(5753) <= data_in(3507);
     data_out(5754) <= data_in(3511);
     data_out(5755) <= data_in(3512);
     data_out(5756) <= data_in(3514);
     data_out(5757) <= data_in(3518);
     data_out(5758) <= data_in(3519);
     data_out(5759) <= data_in(3522);
     data_out(5760) <= data_in(3526);
     data_out(5761) <= data_in(3529);
     data_out(5762) <= data_in(3534);
     data_out(5763) <= data_in(3536);
     data_out(5764) <= data_in(3537);
     data_out(5765) <= data_in(3539);
     data_out(5766) <= data_in(3540);
     data_out(5767) <= data_in(3541);
     data_out(5768) <= data_in(3542);
     data_out(5769) <= data_in(3543);
     data_out(5770) <= data_in(3547);
     data_out(5771) <= data_in(3548);
     data_out(5772) <= data_in(3549);
     data_out(5773) <= data_in(3554);
     data_out(5774) <= data_in(3555);
     data_out(5775) <= data_in(3558);
     data_out(5776) <= data_in(3559);
     data_out(5777) <= data_in(3562);
     data_out(5778) <= data_in(3563);
     data_out(5779) <= data_in(3565);
     data_out(5780) <= data_in(3567);
     data_out(5781) <= data_in(3572);
     data_out(5782) <= data_in(3573);
     data_out(5783) <= data_in(3578);
     data_out(5784) <= data_in(3580);
     data_out(5785) <= data_in(3581);
     data_out(5786) <= data_in(3582);
     data_out(5787) <= data_in(3584);
     data_out(5788) <= data_in(3586);
     data_out(5789) <= data_in(3594);
     data_out(5790) <= data_in(3595);
     data_out(5791) <= data_in(3598);
     data_out(5792) <= data_in(3599);
     data_out(5793) <= data_in(3603);
     data_out(5794) <= data_in(3610);
     data_out(5795) <= data_in(3612);
     data_out(5796) <= data_in(3618);
     data_out(5797) <= data_in(3619);
     data_out(5798) <= data_in(3621);
     data_out(5799) <= data_in(3623);
     data_out(5800) <= data_in(3625);
     data_out(5801) <= data_in(3626);
     data_out(5802) <= data_in(3627);
     data_out(5803) <= data_in(3628);
     data_out(5804) <= data_in(3630);
     data_out(5805) <= data_in(3633);
     data_out(5806) <= data_in(3636);
     data_out(5807) <= data_in(3637);
     data_out(5808) <= data_in(3642);
     data_out(5809) <= data_in(3643);
     data_out(5810) <= data_in(3644);
     data_out(5811) <= data_in(3645);
     data_out(5812) <= data_in(3650);
     data_out(5813) <= data_in(3656);
     data_out(5814) <= data_in(3658);
     data_out(5815) <= data_in(3659);
     data_out(5816) <= data_in(3663);
     data_out(5817) <= data_in(3665);
     data_out(5818) <= data_in(3666);
     data_out(5819) <= data_in(3667);
     data_out(5820) <= data_in(3669);
     data_out(5821) <= data_in(3679);
     data_out(5822) <= data_in(3680);
     data_out(5823) <= data_in(3681);
     data_out(5824) <= data_in(3682);
     data_out(5825) <= data_in(3683);
     data_out(5826) <= data_in(3685);
     data_out(5827) <= data_in(3687);
     data_out(5828) <= data_in(3688);
     data_out(5829) <= data_in(3689);
     data_out(5830) <= data_in(3690);
     data_out(5831) <= data_in(3696);
     data_out(5832) <= data_in(3703);
     data_out(5833) <= data_in(3704);
     data_out(5834) <= data_in(3711);
     data_out(5835) <= data_in(3713);
     data_out(5836) <= data_in(3715);
     data_out(5837) <= data_in(3716);
     data_out(5838) <= data_in(3719);
     data_out(5839) <= data_in(3721);
     data_out(5840) <= data_in(3722);
     data_out(5841) <= data_in(3727);
     data_out(5842) <= data_in(3728);
     data_out(5843) <= data_in(3733);
     data_out(5844) <= data_in(3735);
     data_out(5845) <= data_in(3738);
     data_out(5846) <= data_in(3741);
     data_out(5847) <= data_in(3743);
     data_out(5848) <= data_in(3747);
     data_out(5849) <= data_in(3748);
     data_out(5850) <= data_in(3752);
     data_out(5851) <= data_in(3754);
     data_out(5852) <= data_in(3763);
     data_out(5853) <= data_in(3764);
     data_out(5854) <= data_in(3766);
     data_out(5855) <= data_in(3767);
     data_out(5856) <= data_in(3769);
     data_out(5857) <= data_in(3770);
     data_out(5858) <= data_in(3773);
     data_out(5859) <= data_in(3778);
     data_out(5860) <= data_in(3779);
     data_out(5861) <= data_in(3780);
     data_out(5862) <= data_in(3784);
     data_out(5863) <= data_in(3785);
     data_out(5864) <= data_in(3786);
     data_out(5865) <= data_in(3791);
     data_out(5866) <= data_in(3795);
     data_out(5867) <= data_in(3796);
     data_out(5868) <= data_in(3797);
     data_out(5869) <= data_in(3800);
     data_out(5870) <= data_in(3802);
     data_out(5871) <= data_in(3804);
     data_out(5872) <= data_in(3812);
     data_out(5873) <= data_in(3815);
     data_out(5874) <= data_in(3817);
     data_out(5875) <= data_in(3822);
     data_out(5876) <= data_in(3823);
     data_out(5877) <= data_in(3825);
     data_out(5878) <= data_in(3827);
     data_out(5879) <= data_in(3828);
     data_out(5880) <= data_in(3832);
     data_out(5881) <= data_in(3833);
     data_out(5882) <= data_in(3834);
     data_out(5883) <= data_in(3835);
     data_out(5884) <= data_in(3836);
     data_out(5885) <= data_in(3837);
     data_out(5886) <= data_in(3838);
     data_out(5887) <= data_in(3840);
     data_out(5888) <= data_in(3841);
     data_out(5889) <= data_in(3843);
     data_out(5890) <= data_in(3846);
     data_out(5891) <= data_in(3847);
     data_out(5892) <= data_in(3849);
     data_out(5893) <= data_in(3853);
     data_out(5894) <= data_in(3854);
     data_out(5895) <= data_in(3857);
     data_out(5896) <= data_in(3859);
     data_out(5897) <= data_in(3865);
     data_out(5898) <= data_in(3866);
     data_out(5899) <= data_in(3867);
     data_out(5900) <= data_in(3870);
     data_out(5901) <= data_in(3871);
     data_out(5902) <= data_in(3872);
     data_out(5903) <= data_in(3875);
     data_out(5904) <= data_in(3876);
     data_out(5905) <= data_in(3880);
     data_out(5906) <= data_in(3881);
     data_out(5907) <= data_in(3882);
     data_out(5908) <= data_in(3886);
     data_out(5909) <= data_in(3887);
     data_out(5910) <= data_in(3892);
     data_out(5911) <= data_in(3896);
     data_out(5912) <= data_in(3898);
     data_out(5913) <= data_in(3899);
     data_out(5914) <= data_in(3900);
     data_out(5915) <= data_in(3904);
     data_out(5916) <= data_in(3905);
     data_out(5917) <= data_in(3907);
     data_out(5918) <= data_in(3908);
     data_out(5919) <= data_in(3909);
     data_out(5920) <= data_in(3912);
     data_out(5921) <= data_in(3913);
     data_out(5922) <= data_in(3914);
     data_out(5923) <= data_in(3917);
     data_out(5924) <= data_in(3920);
     data_out(5925) <= data_in(3921);
     data_out(5926) <= data_in(3924);
     data_out(5927) <= data_in(3929);
     data_out(5928) <= data_in(3933);
     data_out(5929) <= data_in(3940);
     data_out(5930) <= data_in(3946);
     data_out(5931) <= data_in(3948);
     data_out(5932) <= data_in(3950);
     data_out(5933) <= data_in(3955);
     data_out(5934) <= data_in(3957);
     data_out(5935) <= data_in(3959);
     data_out(5936) <= data_in(3965);
     data_out(5937) <= data_in(3968);
     data_out(5938) <= data_in(3971);
     data_out(5939) <= data_in(3974);
     data_out(5940) <= data_in(3975);
     data_out(5941) <= data_in(3980);
     data_out(5942) <= data_in(3983);
     data_out(5943) <= data_in(3986);
     data_out(5944) <= data_in(3989);
     data_out(5945) <= data_in(3994);
     data_out(5946) <= data_in(3998);
     data_out(5947) <= data_in(3999);
     data_out(5948) <= data_in(4001);
     data_out(5949) <= data_in(4008);
     data_out(5950) <= data_in(4011);
     data_out(5951) <= data_in(4013);
     data_out(5952) <= data_in(4015);
     data_out(5953) <= data_in(4017);
     data_out(5954) <= data_in(4019);
     data_out(5955) <= data_in(4020);
     data_out(5956) <= data_in(4021);
     data_out(5957) <= data_in(4026);
     data_out(5958) <= data_in(4027);
     data_out(5959) <= data_in(4030);
     data_out(5960) <= data_in(4032);
     data_out(5961) <= data_in(4033);
     data_out(5962) <= data_in(4036);
     data_out(5963) <= data_in(4038);
     data_out(5964) <= data_in(4040);
     data_out(5965) <= data_in(4043);
     data_out(5966) <= data_in(4049);
     data_out(5967) <= data_in(4051);
     data_out(5968) <= data_in(4054);
     data_out(5969) <= data_in(4055);
     data_out(5970) <= data_in(4057);
     data_out(5971) <= data_in(4059);
     data_out(5972) <= data_in(4063);
     data_out(5973) <= data_in(4064);
     data_out(5974) <= data_in(4067);
     data_out(5975) <= data_in(4068);
     data_out(5976) <= data_in(4069);
     data_out(5977) <= data_in(4072);
     data_out(5978) <= data_in(4075);
     data_out(5979) <= data_in(4077);
     data_out(5980) <= data_in(4079);
     data_out(5981) <= data_in(4080);
     data_out(5982) <= data_in(4082);
     data_out(5983) <= data_in(4083);
     data_out(5984) <= data_in(4086);
     data_out(5985) <= data_in(4087);
     data_out(5986) <= data_in(4088);
     data_out(5987) <= data_in(4091);
     data_out(5988) <= data_in(4092);
     data_out(5989) <= data_in(4095);
     data_out(5990) <= data_in(4100);
     data_out(5991) <= data_in(4102);
     data_out(5992) <= data_in(4105);
     data_out(5993) <= data_in(4107);
     data_out(5994) <= data_in(4108);
     data_out(5995) <= data_in(4114);
     data_out(5996) <= data_in(4115);
     data_out(5997) <= data_in(4117);
     data_out(5998) <= data_in(4120);
     data_out(5999) <= data_in(4123);
     data_out(6000) <= data_in(4127);
     data_out(6001) <= data_in(4128);
     data_out(6002) <= data_in(4133);
     data_out(6003) <= data_in(4137);
     data_out(6004) <= data_in(4144);
     data_out(6005) <= data_in(4145);
     data_out(6006) <= data_in(4147);
     data_out(6007) <= data_in(4152);
     data_out(6008) <= data_in(4154);
     data_out(6009) <= data_in(4155);
     data_out(6010) <= data_in(4156);
     data_out(6011) <= data_in(4157);
     data_out(6012) <= data_in(4158);
     data_out(6013) <= data_in(4162);
     data_out(6014) <= data_in(4164);
     data_out(6015) <= data_in(4167);
     data_out(6016) <= data_in(4168);
     data_out(6017) <= data_in(4176);
     data_out(6018) <= data_in(4177);
     data_out(6019) <= data_in(4178);
     data_out(6020) <= data_in(4179);
     data_out(6021) <= data_in(4180);
     data_out(6022) <= data_in(4187);
     data_out(6023) <= data_in(4191);
     data_out(6024) <= data_in(4192);
     data_out(6025) <= data_in(4195);
     data_out(6026) <= data_in(4196);
     data_out(6027) <= data_in(4198);
     data_out(6028) <= data_in(4200);
     data_out(6029) <= data_in(4201);
     data_out(6030) <= data_in(4202);
     data_out(6031) <= data_in(4205);
     data_out(6032) <= data_in(4208);
     data_out(6033) <= data_in(4211);
     data_out(6034) <= data_in(4215);
     data_out(6035) <= data_in(4217);
     data_out(6036) <= data_in(4221);
     data_out(6037) <= data_in(4225);
     data_out(6038) <= data_in(4226);
     data_out(6039) <= data_in(4227);
     data_out(6040) <= data_in(4228);
     data_out(6041) <= data_in(4229);
     data_out(6042) <= data_in(4231);
     data_out(6043) <= data_in(4235);
     data_out(6044) <= data_in(4242);
     data_out(6045) <= data_in(4243);
     data_out(6046) <= data_in(4247);
     data_out(6047) <= data_in(4250);
     data_out(6048) <= data_in(4255);
     data_out(6049) <= data_in(4256);
     data_out(6050) <= data_in(4259);
     data_out(6051) <= data_in(4261);
     data_out(6052) <= data_in(4263);
     data_out(6053) <= data_in(4264);
     data_out(6054) <= data_in(4269);
     data_out(6055) <= data_in(4272);
     data_out(6056) <= data_in(4273);
     data_out(6057) <= data_in(4275);
     data_out(6058) <= data_in(4278);
     data_out(6059) <= data_in(4285);
     data_out(6060) <= data_in(4286);
     data_out(6061) <= data_in(4293);
     data_out(6062) <= data_in(4295);
     data_out(6063) <= data_in(4296);
     data_out(6064) <= data_in(4299);
     data_out(6065) <= data_in(4300);
     data_out(6066) <= data_in(4301);
     data_out(6067) <= data_in(4303);
     data_out(6068) <= data_in(4308);
     data_out(6069) <= data_in(4310);
     data_out(6070) <= data_in(4311);
     data_out(6071) <= data_in(4314);
     data_out(6072) <= data_in(4315);
     data_out(6073) <= data_in(4316);
     data_out(6074) <= data_in(4318);
     data_out(6075) <= data_in(4319);
     data_out(6076) <= data_in(4321);
     data_out(6077) <= data_in(4324);
     data_out(6078) <= data_in(4331);
     data_out(6079) <= data_in(4333);
     data_out(6080) <= data_in(4334);
     data_out(6081) <= data_in(4335);
     data_out(6082) <= data_in(4336);
     data_out(6083) <= data_in(4338);
     data_out(6084) <= data_in(4341);
     data_out(6085) <= data_in(4344);
     data_out(6086) <= data_in(4348);
     data_out(6087) <= data_in(4349);
     data_out(6088) <= data_in(4351);
     data_out(6089) <= data_in(4353);
     data_out(6090) <= data_in(4356);
     data_out(6091) <= data_in(4362);
     data_out(6092) <= data_in(4370);
     data_out(6093) <= data_in(4373);
     data_out(6094) <= data_in(4374);
     data_out(6095) <= data_in(4378);
     data_out(6096) <= data_in(4381);
     data_out(6097) <= data_in(4386);
     data_out(6098) <= data_in(4389);
     data_out(6099) <= data_in(4394);
     data_out(6100) <= data_in(4395);
     data_out(6101) <= data_in(4396);
     data_out(6102) <= data_in(4397);
     data_out(6103) <= data_in(4398);
     data_out(6104) <= data_in(4399);
     data_out(6105) <= data_in(4400);
     data_out(6106) <= data_in(4401);
     data_out(6107) <= data_in(4403);
     data_out(6108) <= data_in(4405);
     data_out(6109) <= data_in(4410);
     data_out(6110) <= data_in(4411);
     data_out(6111) <= data_in(4413);
     data_out(6112) <= data_in(4414);
     data_out(6113) <= data_in(4415);
     data_out(6114) <= data_in(4419);
     data_out(6115) <= data_in(4421);
     data_out(6116) <= data_in(4423);
     data_out(6117) <= data_in(4427);
     data_out(6118) <= data_in(4430);
     data_out(6119) <= data_in(4432);
     data_out(6120) <= data_in(4433);
     data_out(6121) <= data_in(4436);
     data_out(6122) <= data_in(4437);
     data_out(6123) <= data_in(4438);
     data_out(6124) <= data_in(4440);
     data_out(6125) <= data_in(4441);
     data_out(6126) <= data_in(4443);
     data_out(6127) <= data_in(4445);
     data_out(6128) <= data_in(4452);
     data_out(6129) <= data_in(4455);
     data_out(6130) <= data_in(4460);
     data_out(6131) <= data_in(4464);
     data_out(6132) <= data_in(4465);
     data_out(6133) <= data_in(4466);
     data_out(6134) <= data_in(4469);
     data_out(6135) <= data_in(4470);
     data_out(6136) <= data_in(4472);
     data_out(6137) <= data_in(4476);
     data_out(6138) <= data_in(4477);
     data_out(6139) <= data_in(4481);
     data_out(6140) <= data_in(4482);
     data_out(6141) <= data_in(4487);
     data_out(6142) <= data_in(4490);
     data_out(6143) <= data_in(4492);
     data_out(6144) <= data_in(4494);
     data_out(6145) <= data_in(4504);
     data_out(6146) <= data_in(4507);
     data_out(6147) <= data_in(4509);
     data_out(6148) <= data_in(4512);
     data_out(6149) <= data_in(4515);
     data_out(6150) <= data_in(4517);
     data_out(6151) <= data_in(4520);
     data_out(6152) <= data_in(4521);
     data_out(6153) <= data_in(4526);
     data_out(6154) <= data_in(4530);
     data_out(6155) <= data_in(4531);
     data_out(6156) <= data_in(4536);
     data_out(6157) <= data_in(4537);
     data_out(6158) <= data_in(4542);
     data_out(6159) <= data_in(4546);
     data_out(6160) <= data_in(4553);
     data_out(6161) <= data_in(4556);
     data_out(6162) <= data_in(4559);
     data_out(6163) <= data_in(4562);
     data_out(6164) <= data_in(4574);
     data_out(6165) <= data_in(4578);
     data_out(6166) <= data_in(4580);
     data_out(6167) <= data_in(4581);
     data_out(6168) <= data_in(4583);
     data_out(6169) <= data_in(4585);
     data_out(6170) <= data_in(4595);
     data_out(6171) <= data_in(4597);
     data_out(6172) <= data_in(4598);
     data_out(6173) <= data_in(4600);
     data_out(6174) <= data_in(4601);
     data_out(6175) <= data_in(4602);
     data_out(6176) <= data_in(4610);
     data_out(6177) <= data_in(4614);
     data_out(6178) <= data_in(4615);
     data_out(6179) <= data_in(4617);
     data_out(6180) <= data_in(4618);
     data_out(6181) <= data_in(4619);
     data_out(6182) <= data_in(4620);
     data_out(6183) <= data_in(4630);
     data_out(6184) <= data_in(4631);
     data_out(6185) <= data_in(4632);
     data_out(6186) <= data_in(4633);
     data_out(6187) <= data_in(4636);
     data_out(6188) <= data_in(4639);
     data_out(6189) <= data_in(4640);
     data_out(6190) <= data_in(4643);
     data_out(6191) <= data_in(4650);
     data_out(6192) <= data_in(4652);
     data_out(6193) <= data_in(4655);
     data_out(6194) <= data_in(4658);
     data_out(6195) <= data_in(4661);
     data_out(6196) <= data_in(4662);
     data_out(6197) <= data_in(4664);
     data_out(6198) <= data_in(4666);
     data_out(6199) <= data_in(4667);
     data_out(6200) <= data_in(4668);
     data_out(6201) <= data_in(4676);
     data_out(6202) <= data_in(4678);
     data_out(6203) <= data_in(4680);
     data_out(6204) <= data_in(4681);
     data_out(6205) <= data_in(4682);
     data_out(6206) <= data_in(4684);
     data_out(6207) <= data_in(4685);
     data_out(6208) <= data_in(4687);
     data_out(6209) <= data_in(4688);
     data_out(6210) <= data_in(4690);
     data_out(6211) <= data_in(4692);
     data_out(6212) <= data_in(4693);
     data_out(6213) <= data_in(4695);
     data_out(6214) <= data_in(4699);
     data_out(6215) <= data_in(4700);
     data_out(6216) <= data_in(4703);
     data_out(6217) <= data_in(4706);
     data_out(6218) <= data_in(4708);
     data_out(6219) <= data_in(4709);
     data_out(6220) <= data_in(4714);
     data_out(6221) <= data_in(4722);
     data_out(6222) <= data_in(4727);
     data_out(6223) <= data_in(4728);
     data_out(6224) <= data_in(4729);
     data_out(6225) <= data_in(4733);
     data_out(6226) <= data_in(4734);
     data_out(6227) <= data_in(4735);
     data_out(6228) <= data_in(4736);
     data_out(6229) <= data_in(4737);
     data_out(6230) <= data_in(4738);
     data_out(6231) <= data_in(4740);
     data_out(6232) <= data_in(4752);
     data_out(6233) <= data_in(4753);
     data_out(6234) <= data_in(4757);
     data_out(6235) <= data_in(4759);
     data_out(6236) <= data_in(4762);
     data_out(6237) <= data_in(4764);
     data_out(6238) <= data_in(4767);
     data_out(6239) <= data_in(4770);
     data_out(6240) <= data_in(4772);
     data_out(6241) <= data_in(4774);
     data_out(6242) <= data_in(4776);
     data_out(6243) <= data_in(4778);
     data_out(6244) <= data_in(4779);
     data_out(6245) <= data_in(4781);
     data_out(6246) <= data_in(4784);
     data_out(6247) <= data_in(4788);
     data_out(6248) <= data_in(4789);
     data_out(6249) <= data_in(4792);
     data_out(6250) <= data_in(4795);
     data_out(6251) <= data_in(4797);
     data_out(6252) <= data_in(4798);
     data_out(6253) <= data_in(4800);
     data_out(6254) <= data_in(4807);
     data_out(6255) <= data_in(4808);
     data_out(6256) <= data_in(4814);
     data_out(6257) <= data_in(4819);
     data_out(6258) <= data_in(4824);
     data_out(6259) <= data_in(4828);
     data_out(6260) <= data_in(4832);
     data_out(6261) <= data_in(4836);
     data_out(6262) <= data_in(4837);
     data_out(6263) <= data_in(4838);
     data_out(6264) <= data_in(4840);
     data_out(6265) <= data_in(4843);
     data_out(6266) <= data_in(4847);
     data_out(6267) <= data_in(4849);
     data_out(6268) <= data_in(4854);
     data_out(6269) <= data_in(4856);
     data_out(6270) <= data_in(4858);
     data_out(6271) <= data_in(4863);
     data_out(6272) <= data_in(4869);
     data_out(6273) <= data_in(4870);
     data_out(6274) <= data_in(4872);
     data_out(6275) <= data_in(4877);
     data_out(6276) <= data_in(4878);
     data_out(6277) <= data_in(4880);
     data_out(6278) <= data_in(4881);
     data_out(6279) <= data_in(4882);
     data_out(6280) <= data_in(4885);
     data_out(6281) <= data_in(4888);
     data_out(6282) <= data_in(4889);
     data_out(6283) <= data_in(4894);
     data_out(6284) <= data_in(4898);
     data_out(6285) <= data_in(4899);
     data_out(6286) <= data_in(4903);
     data_out(6287) <= data_in(4906);
     data_out(6288) <= data_in(4910);
     data_out(6289) <= data_in(4913);
     data_out(6290) <= data_in(4920);
     data_out(6291) <= data_in(4925);
     data_out(6292) <= data_in(4930);
     data_out(6293) <= data_in(4937);
     data_out(6294) <= data_in(4940);
     data_out(6295) <= data_in(4942);
     data_out(6296) <= data_in(4943);
     data_out(6297) <= data_in(4948);
     data_out(6298) <= data_in(4950);
     data_out(6299) <= data_in(4952);
     data_out(6300) <= data_in(4954);
     data_out(6301) <= data_in(4955);
     data_out(6302) <= data_in(4957);
     data_out(6303) <= data_in(4961);
     data_out(6304) <= data_in(4963);
     data_out(6305) <= data_in(4964);
     data_out(6306) <= data_in(4966);
     data_out(6307) <= data_in(4967);
     data_out(6308) <= data_in(4969);
     data_out(6309) <= data_in(4972);
     data_out(6310) <= data_in(4973);
     data_out(6311) <= data_in(4978);
     data_out(6312) <= data_in(4979);
     data_out(6313) <= data_in(4984);
     data_out(6314) <= data_in(4985);
     data_out(6315) <= data_in(4986);
     data_out(6316) <= data_in(4991);
     data_out(6317) <= data_in(4995);
     data_out(6318) <= data_in(4996);
     data_out(6319) <= data_in(5000);
     data_out(6320) <= data_in(5002);
     data_out(6321) <= data_in(5003);
     data_out(6322) <= data_in(5004);
     data_out(6323) <= data_in(5005);
     data_out(6324) <= data_in(5006);
     data_out(6325) <= data_in(5008);
     data_out(6326) <= data_in(5010);
     data_out(6327) <= data_in(5011);
     data_out(6328) <= data_in(5012);
     data_out(6329) <= data_in(5018);
     data_out(6330) <= data_in(5019);
     data_out(6331) <= data_in(5022);
     data_out(6332) <= data_in(5025);
     data_out(6333) <= data_in(5029);
     data_out(6334) <= data_in(5032);
     data_out(6335) <= data_in(5036);
     data_out(6336) <= data_in(5037);
     data_out(6337) <= data_in(5038);
     data_out(6338) <= data_in(5043);
     data_out(6339) <= data_in(5045);
     data_out(6340) <= data_in(5047);
     data_out(6341) <= data_in(5048);
     data_out(6342) <= data_in(5056);
     data_out(6343) <= data_in(5057);
     data_out(6344) <= data_in(5059);
     data_out(6345) <= data_in(5060);
     data_out(6346) <= data_in(5061);
     data_out(6347) <= data_in(5063);
     data_out(6348) <= data_in(5064);
     data_out(6349) <= data_in(5065);
     data_out(6350) <= data_in(5068);
     data_out(6351) <= data_in(5070);
     data_out(6352) <= data_in(5071);
     data_out(6353) <= data_in(5074);
     data_out(6354) <= data_in(5075);
     data_out(6355) <= data_in(5076);
     data_out(6356) <= data_in(5078);
     data_out(6357) <= data_in(5079);
     data_out(6358) <= data_in(5080);
     data_out(6359) <= data_in(5081);
     data_out(6360) <= data_in(5084);
     data_out(6361) <= data_in(5085);
     data_out(6362) <= data_in(5092);
     data_out(6363) <= data_in(5094);
     data_out(6364) <= data_in(5096);
     data_out(6365) <= data_in(5099);
     data_out(6366) <= data_in(5102);
     data_out(6367) <= data_in(5103);
     data_out(6368) <= data_in(5105);
     data_out(6369) <= data_in(5106);
     data_out(6370) <= data_in(5107);
     data_out(6371) <= data_in(5108);
     data_out(6372) <= data_in(5112);
     data_out(6373) <= data_in(5113);
     data_out(6374) <= data_in(5115);
     data_out(6375) <= data_in(5119);
     data_out(6376) <= data_in(5120);
     data_out(6377) <= data_in(5122);
     data_out(6378) <= data_in(5124);
     data_out(6379) <= data_in(5125);
     data_out(6380) <= data_in(5126);
     data_out(6381) <= data_in(5128);
     data_out(6382) <= data_in(5130);
     data_out(6383) <= data_in(5136);
     data_out(6384) <= data_in(5137);
     data_out(6385) <= data_in(5138);
     data_out(6386) <= data_in(5140);
     data_out(6387) <= data_in(5147);
     data_out(6388) <= data_in(5150);
     data_out(6389) <= data_in(5163);
     data_out(6390) <= data_in(5164);
     data_out(6391) <= data_in(5166);
     data_out(6392) <= data_in(5167);
     data_out(6393) <= data_in(5170);
     data_out(6394) <= data_in(5172);
     data_out(6395) <= data_in(5178);
     data_out(6396) <= data_in(5183);
     data_out(6397) <= data_in(5188);
     data_out(6398) <= data_in(5191);
     data_out(6399) <= data_in(5192);
     data_out(6400) <= data_in(5197);
     data_out(6401) <= data_in(5198);
     data_out(6402) <= data_in(5204);
     data_out(6403) <= data_in(5217);
     data_out(6404) <= data_in(5218);
     data_out(6405) <= data_in(5220);
     data_out(6406) <= data_in(5221);
     data_out(6407) <= data_in(5223);
     data_out(6408) <= data_in(5229);
     data_out(6409) <= data_in(5231);
     data_out(6410) <= data_in(5239);
     data_out(6411) <= data_in(5241);
     data_out(6412) <= data_in(5242);
     data_out(6413) <= data_in(5245);
     data_out(6414) <= data_in(5247);
     data_out(6415) <= data_in(5248);
     data_out(6416) <= data_in(5250);
     data_out(6417) <= data_in(5257);
     data_out(6418) <= data_in(5258);
     data_out(6419) <= data_in(5259);
     data_out(6420) <= data_in(5261);
     data_out(6421) <= data_in(5262);
     data_out(6422) <= data_in(5264);
     data_out(6423) <= data_in(5270);
     data_out(6424) <= data_in(5272);
     data_out(6425) <= data_in(5274);
     data_out(6426) <= data_in(5276);
     data_out(6427) <= data_in(5277);
     data_out(6428) <= data_in(5278);
     data_out(6429) <= data_in(5279);
     data_out(6430) <= data_in(5282);
     data_out(6431) <= data_in(5283);
     data_out(6432) <= data_in(5285);
     data_out(6433) <= data_in(5289);
     data_out(6434) <= data_in(5292);
     data_out(6435) <= data_in(5293);
     data_out(6436) <= data_in(5297);
     data_out(6437) <= data_in(5300);
     data_out(6438) <= data_in(5301);
     data_out(6439) <= data_in(5303);
     data_out(6440) <= data_in(5304);
     data_out(6441) <= data_in(5308);
     data_out(6442) <= data_in(5311);
     data_out(6443) <= data_in(5312);
     data_out(6444) <= data_in(5313);
     data_out(6445) <= data_in(5316);
     data_out(6446) <= data_in(5319);
     data_out(6447) <= data_in(5322);
     data_out(6448) <= data_in(5324);
     data_out(6449) <= data_in(5325);
     data_out(6450) <= data_in(5329);
     data_out(6451) <= data_in(5332);
     data_out(6452) <= data_in(5333);
     data_out(6453) <= data_in(5334);
     data_out(6454) <= data_in(5337);
     data_out(6455) <= data_in(5338);
     data_out(6456) <= data_in(5341);
     data_out(6457) <= data_in(5342);
     data_out(6458) <= data_in(5344);
     data_out(6459) <= data_in(5345);
     data_out(6460) <= data_in(5346);
     data_out(6461) <= data_in(5350);
     data_out(6462) <= data_in(5353);
     data_out(6463) <= data_in(5354);
     data_out(6464) <= data_in(5360);
     data_out(6465) <= data_in(5362);
     data_out(6466) <= data_in(5365);
     data_out(6467) <= data_in(5368);
     data_out(6468) <= data_in(5370);
     data_out(6469) <= data_in(5372);
     data_out(6470) <= data_in(5376);
     data_out(6471) <= data_in(5377);
     data_out(6472) <= data_in(5378);
     data_out(6473) <= data_in(5383);
     data_out(6474) <= data_in(5386);
     data_out(6475) <= data_in(5388);
     data_out(6476) <= data_in(5389);
     data_out(6477) <= data_in(5392);
     data_out(6478) <= data_in(5393);
     data_out(6479) <= data_in(5394);
     data_out(6480) <= data_in(5396);
     data_out(6481) <= data_in(5398);
     data_out(6482) <= data_in(5402);
     data_out(6483) <= data_in(5407);
     data_out(6484) <= data_in(5409);
     data_out(6485) <= data_in(5413);
     data_out(6486) <= data_in(5414);
     data_out(6487) <= data_in(5418);
     data_out(6488) <= data_in(5430);
     data_out(6489) <= data_in(5431);
     data_out(6490) <= data_in(5432);
     data_out(6491) <= data_in(5434);
     data_out(6492) <= data_in(5436);
     data_out(6493) <= data_in(5438);
     data_out(6494) <= data_in(5439);
     data_out(6495) <= data_in(5441);
     data_out(6496) <= data_in(5444);
     data_out(6497) <= data_in(5445);
     data_out(6498) <= data_in(5447);
     data_out(6499) <= data_in(5448);
     data_out(6500) <= data_in(5449);
     data_out(6501) <= data_in(5452);
     data_out(6502) <= data_in(5455);
     data_out(6503) <= data_in(5457);
     data_out(6504) <= data_in(5459);
     data_out(6505) <= data_in(5466);
     data_out(6506) <= data_in(5472);
     data_out(6507) <= data_in(5479);
     data_out(6508) <= data_in(5486);
     data_out(6509) <= data_in(5494);
     data_out(6510) <= data_in(5495);
     data_out(6511) <= data_in(5500);
     data_out(6512) <= data_in(5504);
     data_out(6513) <= data_in(5509);
     data_out(6514) <= data_in(5512);
     data_out(6515) <= data_in(5516);
     data_out(6516) <= data_in(5518);
     data_out(6517) <= data_in(5521);
     data_out(6518) <= data_in(5522);
     data_out(6519) <= data_in(5526);
     data_out(6520) <= data_in(5527);
     data_out(6521) <= data_in(5531);
     data_out(6522) <= data_in(5533);
     data_out(6523) <= data_in(5536);
     data_out(6524) <= data_in(5537);
     data_out(6525) <= data_in(5543);
     data_out(6526) <= data_in(5545);
     data_out(6527) <= data_in(5546);
     data_out(6528) <= data_in(5549);
     data_out(6529) <= data_in(5550);
     data_out(6530) <= data_in(5552);
     data_out(6531) <= data_in(5559);
     data_out(6532) <= data_in(5562);
     data_out(6533) <= data_in(5565);
     data_out(6534) <= data_in(5569);
     data_out(6535) <= data_in(5572);
     data_out(6536) <= data_in(5576);
     data_out(6537) <= data_in(5578);
     data_out(6538) <= data_in(5579);
     data_out(6539) <= data_in(5580);
     data_out(6540) <= data_in(5584);
     data_out(6541) <= data_in(5589);
     data_out(6542) <= data_in(5593);
     data_out(6543) <= data_in(5598);
     data_out(6544) <= data_in(5599);
     data_out(6545) <= data_in(5603);
     data_out(6546) <= data_in(5606);
     data_out(6547) <= data_in(5608);
     data_out(6548) <= data_in(5609);
     data_out(6549) <= data_in(5614);
     data_out(6550) <= data_in(5615);
     data_out(6551) <= data_in(5618);
     data_out(6552) <= data_in(5620);
     data_out(6553) <= data_in(5626);
     data_out(6554) <= data_in(5628);
     data_out(6555) <= data_in(5629);
     data_out(6556) <= data_in(5630);
     data_out(6557) <= data_in(5631);
     data_out(6558) <= data_in(5632);
     data_out(6559) <= data_in(5633);
     data_out(6560) <= data_in(5640);
     data_out(6561) <= data_in(5650);
     data_out(6562) <= data_in(5652);
     data_out(6563) <= data_in(5657);
     data_out(6564) <= data_in(5659);
     data_out(6565) <= data_in(5660);
     data_out(6566) <= data_in(5661);
     data_out(6567) <= data_in(5667);
     data_out(6568) <= data_in(5672);
     data_out(6569) <= data_in(5675);
     data_out(6570) <= data_in(5680);
     data_out(6571) <= data_in(5681);
     data_out(6572) <= data_in(5683);
     data_out(6573) <= data_in(5684);
     data_out(6574) <= data_in(5685);
     data_out(6575) <= data_in(5689);
     data_out(6576) <= data_in(5691);
     data_out(6577) <= data_in(5693);
     data_out(6578) <= data_in(5699);
     data_out(6579) <= data_in(5700);
     data_out(6580) <= data_in(5702);
     data_out(6581) <= data_in(5706);
     data_out(6582) <= data_in(5712);
     data_out(6583) <= data_in(5713);
     data_out(6584) <= data_in(5720);
     data_out(6585) <= data_in(5721);
     data_out(6586) <= data_in(5724);
     data_out(6587) <= data_in(5730);
     data_out(6588) <= data_in(5732);
     data_out(6589) <= data_in(5733);
     data_out(6590) <= data_in(5740);
     data_out(6591) <= data_in(5742);
     data_out(6592) <= data_in(5744);
     data_out(6593) <= data_in(5750);
     data_out(6594) <= data_in(5752);
     data_out(6595) <= data_in(5754);
     data_out(6596) <= data_in(5757);
     data_out(6597) <= data_in(5759);
     data_out(6598) <= data_in(5765);
     data_out(6599) <= data_in(5772);
     data_out(6600) <= data_in(5774);
     data_out(6601) <= data_in(5776);
     data_out(6602) <= data_in(5777);
     data_out(6603) <= data_in(5778);
     data_out(6604) <= data_in(5779);
     data_out(6605) <= data_in(5783);
     data_out(6606) <= data_in(5785);
     data_out(6607) <= data_in(5791);
     data_out(6608) <= data_in(5797);
     data_out(6609) <= data_in(5803);
     data_out(6610) <= data_in(5804);
     data_out(6611) <= data_in(5805);
     data_out(6612) <= data_in(5814);
     data_out(6613) <= data_in(5815);
     data_out(6614) <= data_in(5816);
     data_out(6615) <= data_in(5817);
     data_out(6616) <= data_in(5819);
     data_out(6617) <= data_in(5823);
     data_out(6618) <= data_in(5824);
     data_out(6619) <= data_in(5825);
     data_out(6620) <= data_in(5829);
     data_out(6621) <= data_in(5831);
     data_out(6622) <= data_in(5835);
     data_out(6623) <= data_in(5840);
     data_out(6624) <= data_in(5842);
     data_out(6625) <= data_in(5843);
     data_out(6626) <= data_in(5846);
     data_out(6627) <= data_in(5848);
     data_out(6628) <= data_in(5852);
     data_out(6629) <= data_in(5856);
     data_out(6630) <= data_in(5858);
     data_out(6631) <= data_in(5862);
     data_out(6632) <= data_in(5863);
     data_out(6633) <= data_in(5864);
     data_out(6634) <= data_in(5865);
     data_out(6635) <= data_in(5867);
     data_out(6636) <= data_in(5870);
     data_out(6637) <= data_in(5871);
     data_out(6638) <= data_in(5872);
     data_out(6639) <= data_in(5874);
     data_out(6640) <= data_in(5876);
     data_out(6641) <= data_in(5879);
     data_out(6642) <= data_in(5880);
     data_out(6643) <= data_in(5881);
     data_out(6644) <= data_in(5883);
     data_out(6645) <= data_in(5887);
     data_out(6646) <= data_in(5890);
     data_out(6647) <= data_in(5894);
     data_out(6648) <= data_in(5898);
     data_out(6649) <= data_in(5901);
     data_out(6650) <= data_in(5903);
     data_out(6651) <= data_in(5905);
     data_out(6652) <= data_in(5906);
     data_out(6653) <= data_in(5907);
     data_out(6654) <= data_in(5908);
     data_out(6655) <= data_in(5912);
     data_out(6656) <= data_in(5914);
     data_out(6657) <= data_in(5921);
     data_out(6658) <= data_in(5923);
     data_out(6659) <= data_in(5925);
     data_out(6660) <= data_in(5928);
     data_out(6661) <= data_in(5930);
     data_out(6662) <= data_in(5931);
     data_out(6663) <= data_in(5932);
     data_out(6664) <= data_in(5937);
     data_out(6665) <= data_in(5938);
     data_out(6666) <= data_in(5942);
     data_out(6667) <= data_in(5943);
     data_out(6668) <= data_in(5945);
     data_out(6669) <= data_in(5950);
     data_out(6670) <= data_in(5953);
     data_out(6671) <= data_in(5954);
     data_out(6672) <= data_in(5956);
     data_out(6673) <= data_in(5958);
     data_out(6674) <= data_in(5959);
     data_out(6675) <= data_in(5967);
     data_out(6676) <= data_in(5971);
     data_out(6677) <= data_in(5974);
     data_out(6678) <= data_in(5975);
     data_out(6679) <= data_in(5976);
     data_out(6680) <= data_in(5979);
     data_out(6681) <= data_in(5981);
     data_out(6682) <= data_in(5985);
     data_out(6683) <= data_in(5986);
     data_out(6684) <= data_in(5987);
     data_out(6685) <= data_in(5992);
     data_out(6686) <= data_in(5997);
     data_out(6687) <= data_in(5998);
     data_out(6688) <= data_in(5999);
     data_out(6689) <= data_in(6003);
     data_out(6690) <= data_in(6011);
     data_out(6691) <= data_in(6013);
     data_out(6692) <= data_in(6014);
     data_out(6693) <= data_in(6016);
     data_out(6694) <= data_in(6018);
     data_out(6695) <= data_in(6019);
     data_out(6696) <= data_in(6020);
     data_out(6697) <= data_in(6022);
     data_out(6698) <= data_in(6025);
     data_out(6699) <= data_in(6029);
     data_out(6700) <= data_in(6034);
     data_out(6701) <= data_in(6035);
     data_out(6702) <= data_in(6039);
     data_out(6703) <= data_in(6043);
     data_out(6704) <= data_in(6046);
     data_out(6705) <= data_in(6047);
     data_out(6706) <= data_in(6052);
     data_out(6707) <= data_in(6053);
     data_out(6708) <= data_in(6057);
     data_out(6709) <= data_in(6059);
     data_out(6710) <= data_in(6060);
     data_out(6711) <= data_in(6065);
     data_out(6712) <= data_in(6069);
     data_out(6713) <= data_in(6072);
     data_out(6714) <= data_in(6073);
     data_out(6715) <= data_in(6076);
     data_out(6716) <= data_in(6080);
     data_out(6717) <= data_in(6082);
     data_out(6718) <= data_in(6083);
     data_out(6719) <= data_in(6084);
     data_out(6720) <= data_in(6087);
     data_out(6721) <= data_in(6089);
     data_out(6722) <= data_in(6093);
     data_out(6723) <= data_in(6094);
     data_out(6724) <= data_in(6095);
     data_out(6725) <= data_in(6098);
     data_out(6726) <= data_in(6101);
     data_out(6727) <= data_in(6103);
     data_out(6728) <= data_in(6104);
     data_out(6729) <= data_in(6105);
     data_out(6730) <= data_in(6113);
     data_out(6731) <= data_in(6114);
     data_out(6732) <= data_in(6118);
     data_out(6733) <= data_in(6121);
     data_out(6734) <= data_in(6125);
     data_out(6735) <= data_in(6133);
     data_out(6736) <= data_in(6134);
     data_out(6737) <= data_in(6135);
     data_out(6738) <= data_in(6141);
     data_out(6739) <= data_in(6142);
     data_out(6740) <= data_in(6143);
     data_out(6741) <= data_in(6146);
     data_out(6742) <= data_in(6147);
     data_out(6743) <= data_in(6149);
     data_out(6744) <= data_in(6155);
     data_out(6745) <= data_in(6156);
     data_out(6746) <= data_in(6159);
     data_out(6747) <= data_in(6163);
     data_out(6748) <= data_in(6165);
     data_out(6749) <= data_in(6169);
     data_out(6750) <= data_in(6174);
     data_out(6751) <= data_in(6177);
     data_out(6752) <= data_in(6180);
     data_out(6753) <= data_in(6183);
     data_out(6754) <= data_in(6187);
     data_out(6755) <= data_in(6188);
     data_out(6756) <= data_in(6189);
     data_out(6757) <= data_in(6190);
     data_out(6758) <= data_in(6191);
     data_out(6759) <= data_in(6193);
     data_out(6760) <= data_in(6195);
     data_out(6761) <= data_in(6196);
     data_out(6762) <= data_in(6199);
     data_out(6763) <= data_in(6200);
     data_out(6764) <= data_in(6202);
     data_out(6765) <= data_in(6203);
     data_out(6766) <= data_in(6205);
     data_out(6767) <= data_in(6211);
     data_out(6768) <= data_in(6212);
     data_out(6769) <= data_in(6213);
     data_out(6770) <= data_in(6219);
     data_out(6771) <= data_in(6222);
     data_out(6772) <= data_in(6224);
     data_out(6773) <= data_in(6227);
     data_out(6774) <= data_in(6228);
     data_out(6775) <= data_in(6229);
     data_out(6776) <= data_in(6232);
     data_out(6777) <= data_in(6233);
     data_out(6778) <= data_in(6240);
     data_out(6779) <= data_in(6241);
     data_out(6780) <= data_in(6243);
     data_out(6781) <= data_in(6245);
     data_out(6782) <= data_in(6247);
     data_out(6783) <= data_in(6248);
     data_out(6784) <= data_in(6254);
     data_out(6785) <= data_in(6257);
     data_out(6786) <= data_in(6258);
     data_out(6787) <= data_in(6259);
     data_out(6788) <= data_in(6260);
     data_out(6789) <= data_in(6262);
     data_out(6790) <= data_in(6267);
     data_out(6791) <= data_in(6268);
     data_out(6792) <= data_in(6270);
     data_out(6793) <= data_in(6272);
     data_out(6794) <= data_in(6277);
     data_out(6795) <= data_in(6279);
     data_out(6796) <= data_in(6281);
     data_out(6797) <= data_in(6283);
     data_out(6798) <= data_in(6285);
     data_out(6799) <= data_in(6287);
     data_out(6800) <= data_in(6288);
     data_out(6801) <= data_in(6290);
     data_out(6802) <= data_in(6297);
     data_out(6803) <= data_in(6298);
     data_out(6804) <= data_in(6300);
     data_out(6805) <= data_in(6304);
     data_out(6806) <= data_in(6311);
     data_out(6807) <= data_in(6313);
     data_out(6808) <= data_in(6314);
     data_out(6809) <= data_in(6317);
     data_out(6810) <= data_in(6318);
     data_out(6811) <= data_in(6319);
     data_out(6812) <= data_in(6323);
     data_out(6813) <= data_in(6329);
     data_out(6814) <= data_in(6332);
     data_out(6815) <= data_in(6333);
     data_out(6816) <= data_in(6334);
     data_out(6817) <= data_in(6336);
     data_out(6818) <= data_in(6339);
     data_out(6819) <= data_in(6340);
     data_out(6820) <= data_in(6352);
     data_out(6821) <= data_in(6353);
     data_out(6822) <= data_in(6359);
     data_out(6823) <= data_in(6360);
     data_out(6824) <= data_in(6364);
     data_out(6825) <= data_in(6369);
     data_out(6826) <= data_in(6371);
     data_out(6827) <= data_in(6372);
     data_out(6828) <= data_in(6373);
     data_out(6829) <= data_in(6375);
     data_out(6830) <= data_in(6376);
     data_out(6831) <= data_in(6377);
     data_out(6832) <= data_in(6382);
     data_out(6833) <= data_in(6383);
     data_out(6834) <= data_in(6395);
     data_out(6835) <= data_in(6396);
     data_out(6836) <= data_in(6397);
     data_out(6837) <= data_in(6405);
     data_out(6838) <= data_in(6407);
     data_out(6839) <= data_in(6408);
     data_out(6840) <= data_in(6409);
     data_out(6841) <= data_in(6411);
     data_out(6842) <= data_in(6413);
     data_out(6843) <= data_in(6414);
     data_out(6844) <= data_in(6415);
     data_out(6845) <= data_in(6417);
     data_out(6846) <= data_in(6419);
     data_out(6847) <= data_in(6420);
     data_out(6848) <= data_in(6421);
     data_out(6849) <= data_in(6423);
     data_out(6850) <= data_in(6425);
     data_out(6851) <= data_in(6427);
     data_out(6852) <= data_in(6428);
     data_out(6853) <= data_in(6429);
     data_out(6854) <= data_in(6431);
     data_out(6855) <= data_in(6433);
     data_out(6856) <= data_in(6436);
     data_out(6857) <= data_in(6437);
     data_out(6858) <= data_in(6440);
     data_out(6859) <= data_in(6441);
     data_out(6860) <= data_in(6447);
     data_out(6861) <= data_in(6448);
     data_out(6862) <= data_in(6454);
     data_out(6863) <= data_in(6455);
     data_out(6864) <= data_in(6458);
     data_out(6865) <= data_in(6459);
     data_out(6866) <= data_in(6465);
     data_out(6867) <= data_in(6467);
     data_out(6868) <= data_in(6471);
     data_out(6869) <= data_in(6475);
     data_out(6870) <= data_in(6476);
     data_out(6871) <= data_in(6477);
     data_out(6872) <= data_in(6478);
     data_out(6873) <= data_in(6479);
     data_out(6874) <= data_in(6480);
     data_out(6875) <= data_in(6487);
     data_out(6876) <= data_in(6498);
     data_out(6877) <= data_in(6501);
     data_out(6878) <= data_in(6502);
     data_out(6879) <= data_in(6503);
     data_out(6880) <= data_in(6506);
     data_out(6881) <= data_in(6507);
     data_out(6882) <= data_in(6508);
     data_out(6883) <= data_in(6512);
     data_out(6884) <= data_in(6516);
     data_out(6885) <= data_in(6520);
     data_out(6886) <= data_in(6525);
     data_out(6887) <= data_in(6530);
     data_out(6888) <= data_in(6534);
     data_out(6889) <= data_in(6535);
     data_out(6890) <= data_in(6543);
     data_out(6891) <= data_in(6544);
     data_out(6892) <= data_in(6546);
     data_out(6893) <= data_in(6548);
     data_out(6894) <= data_in(6549);
     data_out(6895) <= data_in(6551);
     data_out(6896) <= data_in(6564);
     data_out(6897) <= data_in(6565);
     data_out(6898) <= data_in(6566);
     data_out(6899) <= data_in(6570);
     data_out(6900) <= data_in(6572);
     data_out(6901) <= data_in(6573);
     data_out(6902) <= data_in(6577);
     data_out(6903) <= data_in(6578);
     data_out(6904) <= data_in(6583);
     data_out(6905) <= data_in(6585);
     data_out(6906) <= data_in(6587);
     data_out(6907) <= data_in(6592);
     data_out(6908) <= data_in(6593);
     data_out(6909) <= data_in(6595);
     data_out(6910) <= data_in(6596);
     data_out(6911) <= data_in(6597);
     data_out(6912) <= data_in(6600);
     data_out(6913) <= data_in(6615);
     data_out(6914) <= data_in(6617);
     data_out(6915) <= data_in(6618);
     data_out(6916) <= data_in(6621);
     data_out(6917) <= data_in(6622);
     data_out(6918) <= data_in(6627);
     data_out(6919) <= data_in(6630);
     data_out(6920) <= data_in(6631);
     data_out(6921) <= data_in(6632);
     data_out(6922) <= data_in(6633);
     data_out(6923) <= data_in(6636);
     data_out(6924) <= data_in(6637);
     data_out(6925) <= data_in(6640);
     data_out(6926) <= data_in(6644);
     data_out(6927) <= data_in(6645);
     data_out(6928) <= data_in(6646);
     data_out(6929) <= data_in(6647);
     data_out(6930) <= data_in(6655);
     data_out(6931) <= data_in(6656);
     data_out(6932) <= data_in(6659);
     data_out(6933) <= data_in(6663);
     data_out(6934) <= data_in(6664);
     data_out(6935) <= data_in(6666);
     data_out(6936) <= data_in(6667);
     data_out(6937) <= data_in(6669);
     data_out(6938) <= data_in(6672);
     data_out(6939) <= data_in(6674);
     data_out(6940) <= data_in(6676);
     data_out(6941) <= data_in(6678);
     data_out(6942) <= data_in(6682);
     data_out(6943) <= data_in(6687);
     data_out(6944) <= data_in(6688);
     data_out(6945) <= data_in(6689);
     data_out(6946) <= data_in(6690);
     data_out(6947) <= data_in(6697);
     data_out(6948) <= data_in(6700);
     data_out(6949) <= data_in(6701);
     data_out(6950) <= data_in(6712);
     data_out(6951) <= data_in(6714);
     data_out(6952) <= data_in(6715);
     data_out(6953) <= data_in(6717);
     data_out(6954) <= data_in(6718);
     data_out(6955) <= data_in(6721);
     data_out(6956) <= data_in(6722);
     data_out(6957) <= data_in(6725);
     data_out(6958) <= data_in(6731);
     data_out(6959) <= data_in(6733);
     data_out(6960) <= data_in(6735);
     data_out(6961) <= data_in(6737);
     data_out(6962) <= data_in(6739);
     data_out(6963) <= data_in(6747);
     data_out(6964) <= data_in(6750);
     data_out(6965) <= data_in(6754);
     data_out(6966) <= data_in(6756);
     data_out(6967) <= data_in(6758);
     data_out(6968) <= data_in(6759);
     data_out(6969) <= data_in(6764);
     data_out(6970) <= data_in(6765);
     data_out(6971) <= data_in(6766);
     data_out(6972) <= data_in(6767);
     data_out(6973) <= data_in(6770);
     data_out(6974) <= data_in(6771);
     data_out(6975) <= data_in(6772);
     data_out(6976) <= data_in(6776);
     data_out(6977) <= data_in(6778);
     data_out(6978) <= data_in(6783);
     data_out(6979) <= data_in(6784);
     data_out(6980) <= data_in(6798);
     data_out(6981) <= data_in(6799);
     data_out(6982) <= data_in(6800);
     data_out(6983) <= data_in(6801);
     data_out(6984) <= data_in(6802);
     data_out(6985) <= data_in(6803);
     data_out(6986) <= data_in(6808);
     data_out(6987) <= data_in(6811);
     data_out(6988) <= data_in(6814);
     data_out(6989) <= data_in(6815);
     data_out(6990) <= data_in(6816);
     data_out(6991) <= data_in(6819);
     data_out(6992) <= data_in(6824);
     data_out(6993) <= data_in(6828);
     data_out(6994) <= data_in(6829);
     data_out(6995) <= data_in(6830);
     data_out(6996) <= data_in(6832);
     data_out(6997) <= data_in(6837);
     data_out(6998) <= data_in(6847);
     data_out(6999) <= data_in(6850);
     data_out(7000) <= data_in(6852);
     data_out(7001) <= data_in(6854);
     data_out(7002) <= data_in(6856);
     data_out(7003) <= data_in(6860);
     data_out(7004) <= data_in(6861);
     data_out(7005) <= data_in(6866);
     data_out(7006) <= data_in(6874);
     data_out(7007) <= data_in(6876);
     data_out(7008) <= data_in(6877);
     data_out(7009) <= data_in(6878);
     data_out(7010) <= data_in(6884);
     data_out(7011) <= data_in(6887);
     data_out(7012) <= data_in(6891);
     data_out(7013) <= data_in(6893);
     data_out(7014) <= data_in(6898);
     data_out(7015) <= data_in(6899);
     data_out(7016) <= data_in(6900);
     data_out(7017) <= data_in(6903);
     data_out(7018) <= data_in(6906);
     data_out(7019) <= data_in(6908);
     data_out(7020) <= data_in(6910);
     data_out(7021) <= data_in(6916);
     data_out(7022) <= data_in(6919);
     data_out(7023) <= data_in(6921);
     data_out(7024) <= data_in(6932);
     data_out(7025) <= data_in(6935);
     data_out(7026) <= data_in(6936);
     data_out(7027) <= data_in(6938);
     data_out(7028) <= data_in(6940);
     data_out(7029) <= data_in(6945);
     data_out(7030) <= data_in(6948);
     data_out(7031) <= data_in(6951);
     data_out(7032) <= data_in(6954);
     data_out(7033) <= data_in(6955);
     data_out(7034) <= data_in(6963);
     data_out(7035) <= data_in(6964);
     data_out(7036) <= data_in(6966);
     data_out(7037) <= data_in(6968);
     data_out(7038) <= data_in(6977);
     data_out(7039) <= data_in(6983);
     data_out(7040) <= data_in(6985);
     data_out(7041) <= data_in(6987);
     data_out(7042) <= data_in(6988);
     data_out(7043) <= data_in(6991);
     data_out(7044) <= data_in(6993);
     data_out(7045) <= data_in(6994);
     data_out(7046) <= data_in(6995);
     data_out(7047) <= data_in(6998);
     data_out(7048) <= data_in(6999);
     data_out(7049) <= data_in(7000);
     data_out(7050) <= data_in(7001);
     data_out(7051) <= data_in(7004);
     data_out(7052) <= data_in(7005);
     data_out(7053) <= data_in(7007);
     data_out(7054) <= data_in(7009);
     data_out(7055) <= data_in(7011);
     data_out(7056) <= data_in(7013);
     data_out(7057) <= data_in(7014);
     data_out(7058) <= data_in(7020);
     data_out(7059) <= data_in(7021);
     data_out(7060) <= data_in(7033);
     data_out(7061) <= data_in(7034);
     data_out(7062) <= data_in(7037);
     data_out(7063) <= data_in(7050);
     data_out(7064) <= data_in(7052);
     data_out(7065) <= data_in(7054);
     data_out(7066) <= data_in(7055);
     data_out(7067) <= data_in(7056);
     data_out(7068) <= data_in(7059);
     data_out(7069) <= data_in(7061);
     data_out(7070) <= data_in(7062);
     data_out(7071) <= data_in(7063);
     data_out(7072) <= data_in(7066);
     data_out(7073) <= data_in(7067);
     data_out(7074) <= data_in(7069);
     data_out(7075) <= data_in(7071);
     data_out(7076) <= data_in(7072);
     data_out(7077) <= data_in(7075);
     data_out(7078) <= data_in(7076);
     data_out(7079) <= data_in(7078);
     data_out(7080) <= data_in(7079);
     data_out(7081) <= data_in(7084);
     data_out(7082) <= data_in(7085);
     data_out(7083) <= data_in(7087);
     data_out(7084) <= data_in(7088);
     data_out(7085) <= data_in(7090);
     data_out(7086) <= data_in(7092);
     data_out(7087) <= data_in(7093);
     data_out(7088) <= data_in(7095);
     data_out(7089) <= data_in(7098);
     data_out(7090) <= data_in(7103);
     data_out(7091) <= data_in(7105);
     data_out(7092) <= data_in(7115);
     data_out(7093) <= data_in(7119);
     data_out(7094) <= data_in(7125);
     data_out(7095) <= data_in(7130);
     data_out(7096) <= data_in(7131);
     data_out(7097) <= data_in(7132);
     data_out(7098) <= data_in(7136);
     data_out(7099) <= data_in(7141);
     data_out(7100) <= data_in(7145);
     data_out(7101) <= data_in(7153);
     data_out(7102) <= data_in(7156);
     data_out(7103) <= data_in(7160);
     data_out(7104) <= data_in(7163);
     data_out(7105) <= data_in(7166);
     data_out(7106) <= data_in(7167);
     data_out(7107) <= data_in(7168);
     data_out(7108) <= data_in(7170);
     data_out(7109) <= data_in(7172);
     data_out(7110) <= data_in(7174);
     data_out(7111) <= data_in(7175);
     data_out(7112) <= data_in(7183);
     data_out(7113) <= data_in(7184);
     data_out(7114) <= data_in(7188);
     data_out(7115) <= data_in(7191);
     data_out(7116) <= data_in(7192);
     data_out(7117) <= data_in(7196);
     data_out(7118) <= data_in(7199);
     data_out(7119) <= data_in(7201);
     data_out(7120) <= data_in(7207);
     data_out(7121) <= data_in(7208);
     data_out(7122) <= data_in(7209);
     data_out(7123) <= data_in(7216);
     data_out(7124) <= data_in(7217);
     data_out(7125) <= data_in(7229);
     data_out(7126) <= data_in(7232);
     data_out(7127) <= data_in(7235);
     data_out(7128) <= data_in(7237);
     data_out(7129) <= data_in(7238);
     data_out(7130) <= data_in(7239);
     data_out(7131) <= data_in(7241);
     data_out(7132) <= data_in(7242);
     data_out(7133) <= data_in(7243);
     data_out(7134) <= data_in(7247);
     data_out(7135) <= data_in(7252);
     data_out(7136) <= data_in(7253);
     data_out(7137) <= data_in(7254);
     data_out(7138) <= data_in(7255);
     data_out(7139) <= data_in(7258);
     data_out(7140) <= data_in(7261);
     data_out(7141) <= data_in(7263);
     data_out(7142) <= data_in(7265);
     data_out(7143) <= data_in(7266);
     data_out(7144) <= data_in(7267);
     data_out(7145) <= data_in(7268);
     data_out(7146) <= data_in(7271);
     data_out(7147) <= data_in(7274);
     data_out(7148) <= data_in(7278);
     data_out(7149) <= data_in(7279);
     data_out(7150) <= data_in(7280);
     data_out(7151) <= data_in(7282);
     data_out(7152) <= data_in(7284);
     data_out(7153) <= data_in(7286);
     data_out(7154) <= data_in(7287);
     data_out(7155) <= data_in(7288);
     data_out(7156) <= data_in(7289);
     data_out(7157) <= data_in(7293);
     data_out(7158) <= data_in(7294);
     data_out(7159) <= data_in(7295);
     data_out(7160) <= data_in(7302);
     data_out(7161) <= data_in(7305);
     data_out(7162) <= data_in(7306);
     data_out(7163) <= data_in(7313);
     data_out(7164) <= data_in(7318);
     data_out(7165) <= data_in(7319);
     data_out(7166) <= data_in(7320);
     data_out(7167) <= data_in(7323);
     data_out(7168) <= data_in(7325);
     data_out(7169) <= data_in(7326);
     data_out(7170) <= data_in(7328);
     data_out(7171) <= data_in(7329);
     data_out(7172) <= data_in(7331);
     data_out(7173) <= data_in(7332);
     data_out(7174) <= data_in(7337);
     data_out(7175) <= data_in(7339);
     data_out(7176) <= data_in(7340);
     data_out(7177) <= data_in(7341);
     data_out(7178) <= data_in(7348);
     data_out(7179) <= data_in(7353);
     data_out(7180) <= data_in(7355);
     data_out(7181) <= data_in(7358);
     data_out(7182) <= data_in(7362);
     data_out(7183) <= data_in(7364);
     data_out(7184) <= data_in(7365);
     data_out(7185) <= data_in(7366);
     data_out(7186) <= data_in(7367);
     data_out(7187) <= data_in(7375);
     data_out(7188) <= data_in(7377);
     data_out(7189) <= data_in(7379);
     data_out(7190) <= data_in(7380);
     data_out(7191) <= data_in(7382);
     data_out(7192) <= data_in(7384);
     data_out(7193) <= data_in(7386);
     data_out(7194) <= data_in(7395);
     data_out(7195) <= data_in(7396);
     data_out(7196) <= data_in(7400);
     data_out(7197) <= data_in(7402);
     data_out(7198) <= data_in(7403);
     data_out(7199) <= data_in(7407);
     data_out(7200) <= data_in(7409);
     data_out(7201) <= data_in(7410);
     data_out(7202) <= data_in(7412);
     data_out(7203) <= data_in(7413);
     data_out(7204) <= data_in(7415);
     data_out(7205) <= data_in(7416);
     data_out(7206) <= data_in(7418);
     data_out(7207) <= data_in(7420);
     data_out(7208) <= data_in(7421);
     data_out(7209) <= data_in(7424);
     data_out(7210) <= data_in(7427);
     data_out(7211) <= data_in(7428);
     data_out(7212) <= data_in(7429);
     data_out(7213) <= data_in(7430);
     data_out(7214) <= data_in(7431);
     data_out(7215) <= data_in(7434);
     data_out(7216) <= data_in(7437);
     data_out(7217) <= data_in(7440);
     data_out(7218) <= data_in(7445);
     data_out(7219) <= data_in(7447);
     data_out(7220) <= data_in(7448);
     data_out(7221) <= data_in(7449);
     data_out(7222) <= data_in(7453);
     data_out(7223) <= data_in(7456);
     data_out(7224) <= data_in(7457);
     data_out(7225) <= data_in(7458);
     data_out(7226) <= data_in(7459);
     data_out(7227) <= data_in(7461);
     data_out(7228) <= data_in(7464);
     data_out(7229) <= data_in(7470);
     data_out(7230) <= data_in(7472);
     data_out(7231) <= data_in(7473);
     data_out(7232) <= data_in(7477);
     data_out(7233) <= data_in(7482);
     data_out(7234) <= data_in(7485);
     data_out(7235) <= data_in(7486);
     data_out(7236) <= data_in(7488);
     data_out(7237) <= data_in(7490);
     data_out(7238) <= data_in(7492);
     data_out(7239) <= data_in(7497);
     data_out(7240) <= data_in(7505);
     data_out(7241) <= data_in(7506);
     data_out(7242) <= data_in(7507);
     data_out(7243) <= data_in(7508);
     data_out(7244) <= data_in(7510);
     data_out(7245) <= data_in(7513);
     data_out(7246) <= data_in(7514);
     data_out(7247) <= data_in(7515);
     data_out(7248) <= data_in(7518);
     data_out(7249) <= data_in(7522);
     data_out(7250) <= data_in(7523);
     data_out(7251) <= data_in(7524);
     data_out(7252) <= data_in(7529);
     data_out(7253) <= data_in(7532);
     data_out(7254) <= data_in(7533);
     data_out(7255) <= data_in(7536);
     data_out(7256) <= data_in(7538);
     data_out(7257) <= data_in(7544);
     data_out(7258) <= data_in(7545);
     data_out(7259) <= data_in(7546);
     data_out(7260) <= data_in(7550);
     data_out(7261) <= data_in(7553);
     data_out(7262) <= data_in(7555);
     data_out(7263) <= data_in(7556);
     data_out(7264) <= data_in(7557);
     data_out(7265) <= data_in(7559);
     data_out(7266) <= data_in(7561);
     data_out(7267) <= data_in(7562);
     data_out(7268) <= data_in(7563);
     data_out(7269) <= data_in(7564);
     data_out(7270) <= data_in(7565);
     data_out(7271) <= data_in(7566);
     data_out(7272) <= data_in(7568);
     data_out(7273) <= data_in(7574);
     data_out(7274) <= data_in(7582);
     data_out(7275) <= data_in(7583);
     data_out(7276) <= data_in(7585);
     data_out(7277) <= data_in(7588);
     data_out(7278) <= data_in(7590);
     data_out(7279) <= data_in(7591);
     data_out(7280) <= data_in(7596);
     data_out(7281) <= data_in(7604);
     data_out(7282) <= data_in(7605);
     data_out(7283) <= data_in(7608);
     data_out(7284) <= data_in(7611);
     data_out(7285) <= data_in(7616);
     data_out(7286) <= data_in(7618);
     data_out(7287) <= data_in(7619);
     data_out(7288) <= data_in(7627);
     data_out(7289) <= data_in(7628);
     data_out(7290) <= data_in(7629);
     data_out(7291) <= data_in(7631);
     data_out(7292) <= data_in(7632);
     data_out(7293) <= data_in(7634);
     data_out(7294) <= data_in(7635);
     data_out(7295) <= data_in(7636);
     data_out(7296) <= data_in(7637);
     data_out(7297) <= data_in(7640);
     data_out(7298) <= data_in(7641);
     data_out(7299) <= data_in(7642);
     data_out(7300) <= data_in(7649);
     data_out(7301) <= data_in(7651);
     data_out(7302) <= data_in(7652);
     data_out(7303) <= data_in(7653);
     data_out(7304) <= data_in(7655);
     data_out(7305) <= data_in(7658);
     data_out(7306) <= data_in(7659);
     data_out(7307) <= data_in(7662);
     data_out(7308) <= data_in(7664);
     data_out(7309) <= data_in(7665);
     data_out(7310) <= data_in(7668);
     data_out(7311) <= data_in(7670);
     data_out(7312) <= data_in(7671);
     data_out(7313) <= data_in(7673);
     data_out(7314) <= data_in(7674);
     data_out(7315) <= data_in(7675);
     data_out(7316) <= data_in(7682);
     data_out(7317) <= data_in(7684);
     data_out(7318) <= data_in(7687);
     data_out(7319) <= data_in(7689);
     data_out(7320) <= data_in(7691);
     data_out(7321) <= data_in(7696);
     data_out(7322) <= data_in(7697);
     data_out(7323) <= data_in(7703);
     data_out(7324) <= data_in(7713);
     data_out(7325) <= data_in(7715);
     data_out(7326) <= data_in(7719);
     data_out(7327) <= data_in(7720);
     data_out(7328) <= data_in(7722);
     data_out(7329) <= data_in(7725);
     data_out(7330) <= data_in(7729);
     data_out(7331) <= data_in(7731);
     data_out(7332) <= data_in(7733);
     data_out(7333) <= data_in(7735);
     data_out(7334) <= data_in(7738);
     data_out(7335) <= data_in(7741);
     data_out(7336) <= data_in(7742);
     data_out(7337) <= data_in(7745);
     data_out(7338) <= data_in(7748);
     data_out(7339) <= data_in(7753);
     data_out(7340) <= data_in(7755);
     data_out(7341) <= data_in(7756);
     data_out(7342) <= data_in(7757);
     data_out(7343) <= data_in(7761);
     data_out(7344) <= data_in(7763);
     data_out(7345) <= data_in(7765);
     data_out(7346) <= data_in(7766);
     data_out(7347) <= data_in(7767);
     data_out(7348) <= data_in(7768);
     data_out(7349) <= data_in(7770);
     data_out(7350) <= data_in(7772);
     data_out(7351) <= data_in(7776);
     data_out(7352) <= data_in(7780);
     data_out(7353) <= data_in(7785);
     data_out(7354) <= data_in(7787);
     data_out(7355) <= data_in(7788);
     data_out(7356) <= data_in(7789);
     data_out(7357) <= data_in(7790);
     data_out(7358) <= data_in(7791);
     data_out(7359) <= data_in(7796);
     data_out(7360) <= data_in(7802);
     data_out(7361) <= data_in(7805);
     data_out(7362) <= data_in(7806);
     data_out(7363) <= data_in(7807);
     data_out(7364) <= data_in(7812);
     data_out(7365) <= data_in(7813);
     data_out(7366) <= data_in(7816);
     data_out(7367) <= data_in(7817);
     data_out(7368) <= data_in(7820);
     data_out(7369) <= data_in(7821);
     data_out(7370) <= data_in(7822);
     data_out(7371) <= data_in(7828);
     data_out(7372) <= data_in(7830);
     data_out(7373) <= data_in(7839);
     data_out(7374) <= data_in(7841);
     data_out(7375) <= data_in(7842);
     data_out(7376) <= data_in(7843);
     data_out(7377) <= data_in(7845);
     data_out(7378) <= data_in(7847);
     data_out(7379) <= data_in(7853);
     data_out(7380) <= data_in(7856);
     data_out(7381) <= data_in(7857);
     data_out(7382) <= data_in(7861);
     data_out(7383) <= data_in(7863);
     data_out(7384) <= data_in(7866);
     data_out(7385) <= data_in(7867);
     data_out(7386) <= data_in(7871);
     data_out(7387) <= data_in(7876);
     data_out(7388) <= data_in(7877);
     data_out(7389) <= data_in(7878);
     data_out(7390) <= data_in(7885);
     data_out(7391) <= data_in(7887);
     data_out(7392) <= data_in(7892);
     data_out(7393) <= data_in(7901);
     data_out(7394) <= data_in(7902);
     data_out(7395) <= data_in(7903);
     data_out(7396) <= data_in(7906);
     data_out(7397) <= data_in(7913);
     data_out(7398) <= data_in(7916);
     data_out(7399) <= data_in(7919);
     data_out(7400) <= data_in(7921);
     data_out(7401) <= data_in(7925);
     data_out(7402) <= data_in(7928);
     data_out(7403) <= data_in(7929);
     data_out(7404) <= data_in(7930);
     data_out(7405) <= data_in(7934);
     data_out(7406) <= data_in(7935);
     data_out(7407) <= data_in(7942);
     data_out(7408) <= data_in(7943);
     data_out(7409) <= data_in(7946);
     data_out(7410) <= data_in(7949);
     data_out(7411) <= data_in(7951);
     data_out(7412) <= data_in(7955);
     data_out(7413) <= data_in(7956);
     data_out(7414) <= data_in(7957);
     data_out(7415) <= data_in(7959);
     data_out(7416) <= data_in(7962);
     data_out(7417) <= data_in(7965);
     data_out(7418) <= data_in(7966);
     data_out(7419) <= data_in(7968);
     data_out(7420) <= data_in(7973);
     data_out(7421) <= data_in(7975);
     data_out(7422) <= data_in(7978);
     data_out(7423) <= data_in(7979);
     data_out(7424) <= data_in(7981);
     data_out(7425) <= data_in(7982);
     data_out(7426) <= data_in(7985);
     data_out(7427) <= data_in(7988);
     data_out(7428) <= data_in(7990);
     data_out(7429) <= data_in(7991);
     data_out(7430) <= data_in(7992);
     data_out(7431) <= data_in(7999);
     data_out(7432) <= data_in(8000);
     data_out(7433) <= data_in(8003);
     data_out(7434) <= data_in(8006);
     data_out(7435) <= data_in(8007);
     data_out(7436) <= data_in(8011);
     data_out(7437) <= data_in(8016);
     data_out(7438) <= data_in(8017);
     data_out(7439) <= data_in(8018);
     data_out(7440) <= data_in(8020);
     data_out(7441) <= data_in(8021);
     data_out(7442) <= data_in(8023);
     data_out(7443) <= data_in(8024);
     data_out(7444) <= data_in(8026);
     data_out(7445) <= data_in(8027);
     data_out(7446) <= data_in(8028);
     data_out(7447) <= data_in(8029);
     data_out(7448) <= data_in(8030);
     data_out(7449) <= data_in(8032);
     data_out(7450) <= data_in(8037);
     data_out(7451) <= data_in(8040);
     data_out(7452) <= data_in(8041);
     data_out(7453) <= data_in(8047);
     data_out(7454) <= data_in(8048);
     data_out(7455) <= data_in(8049);
     data_out(7456) <= data_in(8050);
     data_out(7457) <= data_in(8053);
     data_out(7458) <= data_in(8061);
     data_out(7459) <= data_in(8065);
     data_out(7460) <= data_in(8069);
     data_out(7461) <= data_in(8071);
     data_out(7462) <= data_in(8075);
     data_out(7463) <= data_in(8076);
     data_out(7464) <= data_in(8077);
     data_out(7465) <= data_in(8080);
     data_out(7466) <= data_in(8083);
     data_out(7467) <= data_in(8086);
     data_out(7468) <= data_in(8088);
     data_out(7469) <= data_in(8089);
     data_out(7470) <= data_in(8099);
     data_out(7471) <= data_in(8103);
     data_out(7472) <= data_in(8106);
     data_out(7473) <= data_in(8108);
     data_out(7474) <= data_in(8109);
     data_out(7475) <= data_in(8110);
     data_out(7476) <= data_in(8111);
     data_out(7477) <= data_in(8112);
     data_out(7478) <= data_in(8114);
     data_out(7479) <= data_in(8117);
     data_out(7480) <= data_in(8120);
     data_out(7481) <= data_in(8121);
     data_out(7482) <= data_in(8123);
     data_out(7483) <= data_in(8125);
     data_out(7484) <= data_in(8126);
     data_out(7485) <= data_in(8128);
     data_out(7486) <= data_in(8129);
     data_out(7487) <= data_in(8131);
     data_out(7488) <= data_in(8133);
     data_out(7489) <= data_in(8134);
     data_out(7490) <= data_in(8135);
     data_out(7491) <= data_in(8136);
     data_out(7492) <= data_in(8137);
     data_out(7493) <= data_in(8151);
     data_out(7494) <= data_in(8152);
     data_out(7495) <= data_in(8153);
     data_out(7496) <= data_in(8155);
     data_out(7497) <= data_in(8156);
     data_out(7498) <= data_in(8160);
     data_out(7499) <= data_in(8161);
     data_out(7500) <= data_in(8162);
     data_out(7501) <= data_in(8163);
     data_out(7502) <= data_in(8168);
     data_out(7503) <= data_in(8170);
     data_out(7504) <= data_in(8175);
     data_out(7505) <= data_in(8176);
     data_out(7506) <= data_in(8177);
     data_out(7507) <= data_in(8181);
     data_out(7508) <= data_in(8183);
     data_out(7509) <= data_in(8184);
     data_out(7510) <= data_in(8185);
     data_out(7511) <= data_in(8187);
     data_out(7512) <= data_in(8189);
     data_out(7513) <= data_in(8192);
     data_out(7514) <= data_in(8202);
     data_out(7515) <= data_in(8203);
     data_out(7516) <= data_in(8205);
     data_out(7517) <= data_in(8210);
     data_out(7518) <= data_in(8212);
     data_out(7519) <= data_in(8217);
     data_out(7520) <= data_in(8218);
     data_out(7521) <= data_in(8221);
     data_out(7522) <= data_in(8223);
     data_out(7523) <= data_in(8226);
     data_out(7524) <= data_in(8233);
     data_out(7525) <= data_in(8241);
     data_out(7526) <= data_in(8243);
     data_out(7527) <= data_in(8244);
     data_out(7528) <= data_in(8245);
     data_out(7529) <= data_in(8251);
     data_out(7530) <= data_in(8253);
     data_out(7531) <= data_in(8255);
     data_out(7532) <= data_in(8256);
     data_out(7533) <= data_in(8262);
     data_out(7534) <= data_in(8268);
     data_out(7535) <= data_in(8270);
     data_out(7536) <= data_in(8271);
     data_out(7537) <= data_in(8277);
     data_out(7538) <= data_in(8278);
     data_out(7539) <= data_in(8279);
     data_out(7540) <= data_in(8281);
     data_out(7541) <= data_in(8285);
     data_out(7542) <= data_in(8288);
     data_out(7543) <= data_in(8297);
     data_out(7544) <= data_in(8299);
     data_out(7545) <= data_in(8300);
     data_out(7546) <= data_in(8301);
     data_out(7547) <= data_in(8302);
     data_out(7548) <= data_in(8304);
     data_out(7549) <= data_in(8306);
     data_out(7550) <= data_in(8307);
     data_out(7551) <= data_in(8312);
     data_out(7552) <= data_in(8313);
     data_out(7553) <= data_in(8314);
     data_out(7554) <= data_in(8315);
     data_out(7555) <= data_in(8316);
     data_out(7556) <= data_in(8318);
     data_out(7557) <= data_in(8322);
     data_out(7558) <= data_in(8327);
     data_out(7559) <= data_in(8328);
     data_out(7560) <= data_in(8332);
     data_out(7561) <= data_in(8335);
     data_out(7562) <= data_in(8337);
     data_out(7563) <= data_in(8338);
     data_out(7564) <= data_in(8349);
     data_out(7565) <= data_in(8350);
     data_out(7566) <= data_in(8351);
     data_out(7567) <= data_in(8352);
     data_out(7568) <= data_in(8354);
     data_out(7569) <= data_in(8357);
     data_out(7570) <= data_in(8358);
     data_out(7571) <= data_in(8363);
     data_out(7572) <= data_in(8366);
     data_out(7573) <= data_in(8369);
     data_out(7574) <= data_in(8370);
     data_out(7575) <= data_in(8371);
     data_out(7576) <= data_in(8374);
     data_out(7577) <= data_in(8379);
     data_out(7578) <= data_in(8380);
     data_out(7579) <= data_in(8383);
     data_out(7580) <= data_in(8384);
     data_out(7581) <= data_in(8385);
     data_out(7582) <= data_in(8386);
     data_out(7583) <= data_in(8387);
     data_out(7584) <= data_in(8389);
     data_out(7585) <= data_in(8390);
     data_out(7586) <= data_in(8393);
     data_out(7587) <= data_in(8397);
     data_out(7588) <= data_in(8401);
     data_out(7589) <= data_in(8404);
     data_out(7590) <= data_in(8411);
     data_out(7591) <= data_in(8414);
     data_out(7592) <= data_in(8415);
     data_out(7593) <= data_in(8416);
     data_out(7594) <= data_in(8419);
     data_out(7595) <= data_in(8424);
     data_out(7596) <= data_in(8426);
     data_out(7597) <= data_in(8429);
     data_out(7598) <= data_in(8432);
     data_out(7599) <= data_in(8435);
     data_out(7600) <= data_in(8447);
     data_out(7601) <= data_in(8449);
     data_out(7602) <= data_in(8451);
     data_out(7603) <= data_in(8456);
     data_out(7604) <= data_in(8465);
     data_out(7605) <= data_in(8466);
     data_out(7606) <= data_in(8472);
     data_out(7607) <= data_in(8474);
     data_out(7608) <= data_in(8480);
     data_out(7609) <= data_in(8489);
     data_out(7610) <= data_in(8492);
     data_out(7611) <= data_in(8496);
     data_out(7612) <= data_in(8497);
     data_out(7613) <= data_in(8499);
     data_out(7614) <= data_in(8502);
     data_out(7615) <= data_in(8510);
     data_out(7616) <= data_in(8513);
     data_out(7617) <= data_in(8515);
     data_out(7618) <= data_in(8517);
     data_out(7619) <= data_in(8518);
     data_out(7620) <= data_in(8520);
     data_out(7621) <= data_in(8521);
     data_out(7622) <= data_in(8522);
     data_out(7623) <= data_in(8524);
     data_out(7624) <= data_in(8528);
     data_out(7625) <= data_in(8529);
     data_out(7626) <= data_in(8532);
     data_out(7627) <= data_in(8538);
     data_out(7628) <= data_in(8541);
     data_out(7629) <= data_in(8542);
     data_out(7630) <= data_in(8549);
     data_out(7631) <= data_in(8550);
     data_out(7632) <= data_in(8551);
     data_out(7633) <= data_in(8552);
     data_out(7634) <= data_in(8559);
     data_out(7635) <= data_in(8560);
     data_out(7636) <= data_in(8563);
     data_out(7637) <= data_in(8564);
     data_out(7638) <= data_in(8565);
     data_out(7639) <= data_in(8566);
     data_out(7640) <= data_in(8571);
     data_out(7641) <= data_in(8572);
     data_out(7642) <= data_in(8574);
     data_out(7643) <= data_in(8575);
     data_out(7644) <= data_in(8582);
     data_out(7645) <= data_in(8583);
     data_out(7646) <= data_in(8584);
     data_out(7647) <= data_in(8587);
     data_out(7648) <= data_in(8588);
     data_out(7649) <= data_in(8589);
     data_out(7650) <= data_in(8590);
     data_out(7651) <= data_in(8598);
     data_out(7652) <= data_in(8602);
     data_out(7653) <= data_in(8604);
     data_out(7654) <= data_in(8608);
     data_out(7655) <= data_in(8609);
     data_out(7656) <= data_in(8611);
     data_out(7657) <= data_in(8613);
     data_out(7658) <= data_in(8614);
     data_out(7659) <= data_in(8615);
     data_out(7660) <= data_in(8617);
     data_out(7661) <= data_in(8618);
     data_out(7662) <= data_in(8621);
     data_out(7663) <= data_in(8624);
     data_out(7664) <= data_in(8625);
     data_out(7665) <= data_in(8627);
     data_out(7666) <= data_in(8629);
     data_out(7667) <= data_in(8631);
     data_out(7668) <= data_in(8634);
     data_out(7669) <= data_in(8640);
     data_out(7670) <= data_in(8641);
     data_out(7671) <= data_in(8643);
     data_out(7672) <= data_in(8645);
     data_out(7673) <= data_in(8649);
     data_out(7674) <= data_in(8650);
     data_out(7675) <= data_in(8653);
     data_out(7676) <= data_in(8654);
     data_out(7677) <= data_in(8657);
     data_out(7678) <= data_in(8658);
     data_out(7679) <= data_in(8659);
     data_out(7680) <= data_in(8664);
     data_out(7681) <= data_in(8665);
     data_out(7682) <= data_in(8666);
     data_out(7683) <= data_in(8670);
     data_out(7684) <= data_in(8672);
     data_out(7685) <= data_in(8677);
     data_out(7686) <= data_in(8678);
     data_out(7687) <= data_in(8679);
     data_out(7688) <= data_in(8681);
     data_out(7689) <= data_in(8682);
     data_out(7690) <= data_in(8684);
     data_out(7691) <= data_in(8685);
     data_out(7692) <= data_in(8689);
     data_out(7693) <= data_in(8691);
     data_out(7694) <= data_in(8695);
     data_out(7695) <= data_in(8698);
     data_out(7696) <= data_in(8699);
     data_out(7697) <= data_in(8701);
     data_out(7698) <= data_in(8704);
     data_out(7699) <= data_in(8706);
     data_out(7700) <= data_in(8707);
     data_out(7701) <= data_in(8710);
     data_out(7702) <= data_in(8713);
     data_out(7703) <= data_in(8716);
     data_out(7704) <= data_in(8720);
     data_out(7705) <= data_in(8721);
     data_out(7706) <= data_in(8724);
     data_out(7707) <= data_in(8732);
     data_out(7708) <= data_in(8733);
     data_out(7709) <= data_in(8737);
     data_out(7710) <= data_in(8739);
     data_out(7711) <= data_in(8747);
     data_out(7712) <= data_in(8748);
     data_out(7713) <= data_in(8749);
     data_out(7714) <= data_in(8753);
     data_out(7715) <= data_in(8754);
     data_out(7716) <= data_in(8755);
     data_out(7717) <= data_in(8759);
     data_out(7718) <= data_in(8761);
     data_out(7719) <= data_in(8765);
     data_out(7720) <= data_in(8766);
     data_out(7721) <= data_in(8767);
     data_out(7722) <= data_in(8768);
     data_out(7723) <= data_in(8770);
     data_out(7724) <= data_in(8773);
     data_out(7725) <= data_in(8776);
     data_out(7726) <= data_in(8777);
     data_out(7727) <= data_in(8782);
     data_out(7728) <= data_in(8789);
     data_out(7729) <= data_in(8790);
     data_out(7730) <= data_in(8791);
     data_out(7731) <= data_in(8793);
     data_out(7732) <= data_in(8794);
     data_out(7733) <= data_in(8796);
     data_out(7734) <= data_in(8798);
     data_out(7735) <= data_in(8807);
     data_out(7736) <= data_in(8811);
     data_out(7737) <= data_in(8813);
     data_out(7738) <= data_in(8815);
     data_out(7739) <= data_in(8816);
     data_out(7740) <= data_in(8823);
     data_out(7741) <= data_in(8829);
     data_out(7742) <= data_in(8831);
     data_out(7743) <= data_in(8834);
     data_out(7744) <= data_in(8835);
     data_out(7745) <= data_in(8840);
     data_out(7746) <= data_in(8841);
     data_out(7747) <= data_in(8843);
     data_out(7748) <= data_in(8844);
     data_out(7749) <= data_in(8856);
     data_out(7750) <= data_in(8857);
     data_out(7751) <= data_in(8860);
     data_out(7752) <= data_in(8866);
     data_out(7753) <= data_in(8868);
     data_out(7754) <= data_in(8870);
     data_out(7755) <= data_in(8871);
     data_out(7756) <= data_in(8873);
     data_out(7757) <= data_in(8874);
     data_out(7758) <= data_in(8875);
     data_out(7759) <= data_in(8879);
     data_out(7760) <= data_in(8888);
     data_out(7761) <= data_in(8889);
     data_out(7762) <= data_in(8891);
     data_out(7763) <= data_in(8896);
     data_out(7764) <= data_in(8898);
     data_out(7765) <= data_in(8906);
     data_out(7766) <= data_in(8910);
     data_out(7767) <= data_in(8911);
     data_out(7768) <= data_in(8915);
     data_out(7769) <= data_in(8916);
     data_out(7770) <= data_in(8917);
     data_out(7771) <= data_in(8919);
     data_out(7772) <= data_in(8920);
     data_out(7773) <= data_in(8921);
     data_out(7774) <= data_in(8925);
     data_out(7775) <= data_in(8930);
     data_out(7776) <= data_in(8931);
     data_out(7777) <= data_in(8932);
     data_out(7778) <= data_in(8941);
     data_out(7779) <= data_in(8943);
     data_out(7780) <= data_in(8946);
     data_out(7781) <= data_in(8950);
     data_out(7782) <= data_in(8952);
     data_out(7783) <= data_in(8953);
     data_out(7784) <= data_in(8954);
     data_out(7785) <= data_in(8955);
     data_out(7786) <= data_in(8957);
     data_out(7787) <= data_in(8958);
     data_out(7788) <= data_in(8959);
     data_out(7789) <= data_in(8960);
     data_out(7790) <= data_in(8961);
     data_out(7791) <= data_in(8962);
     data_out(7792) <= data_in(8963);
     data_out(7793) <= data_in(8967);
     data_out(7794) <= data_in(8971);
     data_out(7795) <= data_in(8972);
     data_out(7796) <= data_in(8974);
     data_out(7797) <= data_in(8975);
     data_out(7798) <= data_in(8976);
     data_out(7799) <= data_in(8978);
     data_out(7800) <= data_in(8986);
     data_out(7801) <= data_in(8987);
     data_out(7802) <= data_in(8988);
     data_out(7803) <= data_in(8989);
     data_out(7804) <= data_in(8994);
     data_out(7805) <= data_in(8996);
     data_out(7806) <= data_in(8997);
     data_out(7807) <= data_in(9000);
     data_out(7808) <= data_in(9002);
     data_out(7809) <= data_in(9004);
     data_out(7810) <= data_in(9007);
     data_out(7811) <= data_in(9010);
     data_out(7812) <= data_in(9011);
     data_out(7813) <= data_in(9013);
     data_out(7814) <= data_in(9016);
     data_out(7815) <= data_in(9018);
     data_out(7816) <= data_in(9019);
     data_out(7817) <= data_in(9022);
     data_out(7818) <= data_in(9026);
     data_out(7819) <= data_in(9028);
     data_out(7820) <= data_in(9031);
     data_out(7821) <= data_in(9033);
     data_out(7822) <= data_in(9035);
     data_out(7823) <= data_in(9036);
     data_out(7824) <= data_in(9037);
     data_out(7825) <= data_in(9039);
     data_out(7826) <= data_in(9041);
     data_out(7827) <= data_in(9047);
     data_out(7828) <= data_in(9048);
     data_out(7829) <= data_in(9049);
     data_out(7830) <= data_in(9050);
     data_out(7831) <= data_in(9052);
     data_out(7832) <= data_in(9053);
     data_out(7833) <= data_in(9055);
     data_out(7834) <= data_in(9056);
     data_out(7835) <= data_in(9057);
     data_out(7836) <= data_in(9058);
     data_out(7837) <= data_in(9059);
     data_out(7838) <= data_in(9063);
     data_out(7839) <= data_in(9069);
     data_out(7840) <= data_in(9072);
     data_out(7841) <= data_in(9081);
     data_out(7842) <= data_in(9084);
     data_out(7843) <= data_in(9086);
     data_out(7844) <= data_in(9088);
     data_out(7845) <= data_in(9089);
     data_out(7846) <= data_in(9092);
     data_out(7847) <= data_in(9094);
     data_out(7848) <= data_in(9096);
     data_out(7849) <= data_in(9098);
     data_out(7850) <= data_in(9099);
     data_out(7851) <= data_in(9100);
     data_out(7852) <= data_in(9104);
     data_out(7853) <= data_in(9105);
     data_out(7854) <= data_in(9106);
     data_out(7855) <= data_in(9110);
     data_out(7856) <= data_in(9113);
     data_out(7857) <= data_in(9120);
     data_out(7858) <= data_in(9122);
     data_out(7859) <= data_in(9125);
     data_out(7860) <= data_in(9127);
     data_out(7861) <= data_in(9129);
     data_out(7862) <= data_in(9130);
     data_out(7863) <= data_in(9132);
     data_out(7864) <= data_in(9134);
     data_out(7865) <= data_in(9135);
     data_out(7866) <= data_in(9136);
     data_out(7867) <= data_in(9139);
     data_out(7868) <= data_in(9145);
     data_out(7869) <= data_in(9146);
     data_out(7870) <= data_in(9149);
     data_out(7871) <= data_in(9150);
     data_out(7872) <= data_in(9151);
     data_out(7873) <= data_in(9152);
     data_out(7874) <= data_in(9153);
     data_out(7875) <= data_in(9154);
     data_out(7876) <= data_in(9156);
     data_out(7877) <= data_in(9160);
     data_out(7878) <= data_in(9161);
     data_out(7879) <= data_in(9163);
     data_out(7880) <= data_in(9165);
     data_out(7881) <= data_in(9167);
     data_out(7882) <= data_in(9169);
     data_out(7883) <= data_in(9173);
     data_out(7884) <= data_in(9174);
     data_out(7885) <= data_in(9183);
     data_out(7886) <= data_in(9185);
     data_out(7887) <= data_in(9186);
     data_out(7888) <= data_in(9187);
     data_out(7889) <= data_in(9190);
     data_out(7890) <= data_in(9192);
     data_out(7891) <= data_in(9195);
     data_out(7892) <= data_in(9202);
     data_out(7893) <= data_in(9203);
     data_out(7894) <= data_in(9209);
     data_out(7895) <= data_in(9210);
     data_out(7896) <= data_in(9215);
     data_out(7897) <= data_in(9216);
     data_out(7898) <= data_in(9220);
     data_out(7899) <= data_in(9224);
     data_out(7900) <= data_in(9225);
     data_out(7901) <= data_in(9227);
     data_out(7902) <= data_in(9228);
     data_out(7903) <= data_in(9237);
     data_out(7904) <= data_in(9239);
     data_out(7905) <= data_in(9242);
     data_out(7906) <= data_in(9247);
     data_out(7907) <= data_in(9250);
     data_out(7908) <= data_in(9251);
     data_out(7909) <= data_in(9254);
     data_out(7910) <= data_in(9256);
     data_out(7911) <= data_in(9257);
     data_out(7912) <= data_in(9259);
     data_out(7913) <= data_in(9260);
     data_out(7914) <= data_in(9261);
     data_out(7915) <= data_in(9262);
     data_out(7916) <= data_in(9265);
     data_out(7917) <= data_in(9268);
     data_out(7918) <= data_in(9272);
     data_out(7919) <= data_in(9275);
     data_out(7920) <= data_in(9280);
     data_out(7921) <= data_in(9283);
     data_out(7922) <= data_in(9285);
     data_out(7923) <= data_in(9288);
     data_out(7924) <= data_in(9290);
     data_out(7925) <= data_in(9291);
     data_out(7926) <= data_in(9294);
     data_out(7927) <= data_in(9295);
     data_out(7928) <= data_in(9297);
     data_out(7929) <= data_in(9303);
     data_out(7930) <= data_in(9304);
     data_out(7931) <= data_in(9310);
     data_out(7932) <= data_in(9313);
     data_out(7933) <= data_in(9314);
     data_out(7934) <= data_in(9320);
     data_out(7935) <= data_in(9321);
     data_out(7936) <= data_in(9322);
     data_out(7937) <= data_in(9334);
     data_out(7938) <= data_in(9336);
     data_out(7939) <= data_in(9340);
     data_out(7940) <= data_in(9343);
     data_out(7941) <= data_in(9345);
     data_out(7942) <= data_in(9346);
     data_out(7943) <= data_in(9357);
     data_out(7944) <= data_in(9358);
     data_out(7945) <= data_in(9362);
     data_out(7946) <= data_in(9363);
     data_out(7947) <= data_in(9364);
     data_out(7948) <= data_in(9365);
     data_out(7949) <= data_in(9366);
     data_out(7950) <= data_in(9368);
     data_out(7951) <= data_in(9371);
     data_out(7952) <= data_in(9372);
     data_out(7953) <= data_in(9373);
     data_out(7954) <= data_in(9376);
     data_out(7955) <= data_in(9377);
     data_out(7956) <= data_in(9381);
     data_out(7957) <= data_in(9384);
     data_out(7958) <= data_in(9385);
     data_out(7959) <= data_in(9386);
     data_out(7960) <= data_in(9392);
     data_out(7961) <= data_in(9393);
     data_out(7962) <= data_in(9397);
     data_out(7963) <= data_in(9398);
     data_out(7964) <= data_in(9400);
     data_out(7965) <= data_in(9413);
     data_out(7966) <= data_in(9414);
     data_out(7967) <= data_in(9421);
     data_out(7968) <= data_in(9422);
     data_out(7969) <= data_in(9423);
     data_out(7970) <= data_in(9428);
     data_out(7971) <= data_in(9434);
     data_out(7972) <= data_in(9436);
     data_out(7973) <= data_in(9437);
     data_out(7974) <= data_in(9439);
     data_out(7975) <= data_in(9440);
     data_out(7976) <= data_in(9449);
     data_out(7977) <= data_in(9450);
     data_out(7978) <= data_in(9453);
     data_out(7979) <= data_in(9455);
     data_out(7980) <= data_in(9459);
     data_out(7981) <= data_in(9461);
     data_out(7982) <= data_in(9463);
     data_out(7983) <= data_in(9464);
     data_out(7984) <= data_in(9465);
     data_out(7985) <= data_in(9467);
     data_out(7986) <= data_in(9469);
     data_out(7987) <= data_in(9473);
     data_out(7988) <= data_in(9474);
     data_out(7989) <= data_in(9475);
     data_out(7990) <= data_in(9479);
     data_out(7991) <= data_in(9482);
     data_out(7992) <= data_in(9484);
     data_out(7993) <= data_in(9488);
     data_out(7994) <= data_in(9492);
     data_out(7995) <= data_in(9497);
     data_out(7996) <= data_in(9499);
     data_out(7997) <= data_in(9505);
     data_out(7998) <= data_in(9508);
     data_out(7999) <= data_in(9514);
     data_out(8000) <= data_in(9517);
     data_out(8001) <= data_in(9519);
     data_out(8002) <= data_in(9523);
     data_out(8003) <= data_in(9526);
     data_out(8004) <= data_in(9530);
     data_out(8005) <= data_in(9531);
     data_out(8006) <= data_in(9534);
     data_out(8007) <= data_in(9535);
     data_out(8008) <= data_in(9537);
     data_out(8009) <= data_in(9543);
     data_out(8010) <= data_in(9545);
     data_out(8011) <= data_in(9546);
     data_out(8012) <= data_in(9547);
     data_out(8013) <= data_in(9549);
     data_out(8014) <= data_in(9552);
     data_out(8015) <= data_in(9553);
     data_out(8016) <= data_in(9554);
     data_out(8017) <= data_in(9556);
     data_out(8018) <= data_in(9557);
     data_out(8019) <= data_in(9561);
     data_out(8020) <= data_in(9562);
     data_out(8021) <= data_in(9564);
     data_out(8022) <= data_in(9566);
     data_out(8023) <= data_in(9568);
     data_out(8024) <= data_in(9569);
     data_out(8025) <= data_in(9571);
     data_out(8026) <= data_in(9572);
     data_out(8027) <= data_in(9577);
     data_out(8028) <= data_in(9580);
     data_out(8029) <= data_in(9581);
     data_out(8030) <= data_in(9582);
     data_out(8031) <= data_in(9586);
     data_out(8032) <= data_in(9589);
     data_out(8033) <= data_in(9590);
     data_out(8034) <= data_in(9592);
     data_out(8035) <= data_in(9599);
     data_out(8036) <= data_in(9601);
     data_out(8037) <= data_in(9606);
     data_out(8038) <= data_in(9608);
     data_out(8039) <= data_in(9610);
     data_out(8040) <= data_in(9611);
     data_out(8041) <= data_in(9613);
     data_out(8042) <= data_in(9615);
     data_out(8043) <= data_in(9617);
     data_out(8044) <= data_in(9618);
     data_out(8045) <= data_in(9619);
     data_out(8046) <= data_in(9620);
     data_out(8047) <= data_in(9622);
     data_out(8048) <= data_in(9623);
     data_out(8049) <= data_in(9626);
     data_out(8050) <= data_in(9627);
     data_out(8051) <= data_in(9628);
     data_out(8052) <= data_in(9630);
     data_out(8053) <= data_in(9634);
     data_out(8054) <= data_in(9637);
     data_out(8055) <= data_in(9638);
     data_out(8056) <= data_in(9641);
     data_out(8057) <= data_in(9642);
     data_out(8058) <= data_in(9646);
     data_out(8059) <= data_in(9648);
     data_out(8060) <= data_in(9649);
     data_out(8061) <= data_in(9651);
     data_out(8062) <= data_in(9655);
     data_out(8063) <= data_in(9658);
     data_out(8064) <= data_in(9659);
     data_out(8065) <= data_in(9660);
     data_out(8066) <= data_in(9661);
     data_out(8067) <= data_in(9662);
     data_out(8068) <= data_in(9664);
     data_out(8069) <= data_in(9666);
     data_out(8070) <= data_in(9676);
     data_out(8071) <= data_in(9677);
     data_out(8072) <= data_in(9680);
     data_out(8073) <= data_in(9683);
     data_out(8074) <= data_in(9684);
     data_out(8075) <= data_in(9690);
     data_out(8076) <= data_in(9692);
     data_out(8077) <= data_in(9695);
     data_out(8078) <= data_in(9697);
     data_out(8079) <= data_in(9700);
     data_out(8080) <= data_in(9704);
     data_out(8081) <= data_in(9705);
     data_out(8082) <= data_in(9706);
     data_out(8083) <= data_in(9707);
     data_out(8084) <= data_in(9712);
     data_out(8085) <= data_in(9717);
     data_out(8086) <= data_in(9720);
     data_out(8087) <= data_in(9721);
     data_out(8088) <= data_in(9723);
     data_out(8089) <= data_in(9724);
     data_out(8090) <= data_in(9729);
     data_out(8091) <= data_in(9730);
     data_out(8092) <= data_in(9731);
     data_out(8093) <= data_in(9732);
     data_out(8094) <= data_in(9734);
     data_out(8095) <= data_in(9736);
     data_out(8096) <= data_in(9737);
     data_out(8097) <= data_in(9738);
     data_out(8098) <= data_in(9741);
     data_out(8099) <= data_in(9743);
     data_out(8100) <= data_in(9749);
     data_out(8101) <= data_in(9752);
     data_out(8102) <= data_in(9753);
     data_out(8103) <= data_in(9754);
     data_out(8104) <= data_in(9758);
     data_out(8105) <= data_in(9760);
     data_out(8106) <= data_in(9761);
     data_out(8107) <= data_in(9764);
     data_out(8108) <= data_in(9765);
     data_out(8109) <= data_in(9768);
     data_out(8110) <= data_in(9770);
     data_out(8111) <= data_in(9772);
     data_out(8112) <= data_in(9776);
     data_out(8113) <= data_in(9782);
     data_out(8114) <= data_in(9785);
     data_out(8115) <= data_in(9788);
     data_out(8116) <= data_in(9789);
     data_out(8117) <= data_in(9792);
     data_out(8118) <= data_in(9795);
     data_out(8119) <= data_in(9798);
     data_out(8120) <= data_in(9800);
     data_out(8121) <= data_in(9801);
     data_out(8122) <= data_in(9802);
     data_out(8123) <= data_in(9803);
     data_out(8124) <= data_in(9804);
     data_out(8125) <= data_in(9806);
     data_out(8126) <= data_in(9808);
     data_out(8127) <= data_in(9812);
     data_out(8128) <= data_in(9815);
     data_out(8129) <= data_in(9816);
     data_out(8130) <= data_in(9817);
     data_out(8131) <= data_in(9819);
     data_out(8132) <= data_in(9820);
     data_out(8133) <= data_in(9822);
     data_out(8134) <= data_in(9833);
     data_out(8135) <= data_in(9834);
     data_out(8136) <= data_in(9843);
     data_out(8137) <= data_in(9845);
     data_out(8138) <= data_in(9848);
     data_out(8139) <= data_in(9850);
     data_out(8140) <= data_in(9852);
     data_out(8141) <= data_in(9854);
     data_out(8142) <= data_in(9855);
     data_out(8143) <= data_in(9858);
     data_out(8144) <= data_in(9862);
     data_out(8145) <= data_in(9864);
     data_out(8146) <= data_in(9866);
     data_out(8147) <= data_in(9867);
     data_out(8148) <= data_in(9869);
     data_out(8149) <= data_in(9870);
     data_out(8150) <= data_in(9874);
     data_out(8151) <= data_in(9876);
     data_out(8152) <= data_in(9879);
     data_out(8153) <= data_in(9883);
     data_out(8154) <= data_in(9886);
     data_out(8155) <= data_in(9890);
     data_out(8156) <= data_in(9895);
     data_out(8157) <= data_in(9898);
     data_out(8158) <= data_in(9901);
     data_out(8159) <= data_in(9905);
     data_out(8160) <= data_in(9912);
     data_out(8161) <= data_in(9915);
     data_out(8162) <= data_in(9917);
     data_out(8163) <= data_in(9918);
     data_out(8164) <= data_in(9919);
     data_out(8165) <= data_in(9921);
     data_out(8166) <= data_in(9927);
     data_out(8167) <= data_in(9929);
     data_out(8168) <= data_in(9931);
     data_out(8169) <= data_in(9936);
     data_out(8170) <= data_in(9940);
     data_out(8171) <= data_in(9950);
     data_out(8172) <= data_in(9952);
     data_out(8173) <= data_in(9957);
     data_out(8174) <= data_in(9958);
     data_out(8175) <= data_in(9963);
     data_out(8176) <= data_in(9964);
     data_out(8177) <= data_in(9967);
     data_out(8178) <= data_in(9971);
     data_out(8179) <= data_in(9974);
     data_out(8180) <= data_in(9976);
     data_out(8181) <= data_in(9985);
     data_out(8182) <= data_in(9992);
     data_out(8183) <= data_in(9993);
     data_out(8184) <= data_in(9998);
     data_out(8185) <= data_in(10002);
     data_out(8186) <= data_in(10004);
     data_out(8187) <= data_in(10008);
     data_out(8188) <= data_in(10009);
     data_out(8189) <= data_in(10010);
     data_out(8190) <= data_in(10011);
     data_out(8191) <= data_in(10012);
     data_out(8192) <= data_in(10014);
     data_out(8193) <= data_in(10017);
     data_out(8194) <= data_in(10018);
     data_out(8195) <= data_in(10020);
     data_out(8196) <= data_in(10022);
     data_out(8197) <= data_in(10026);
     data_out(8198) <= data_in(10035);
     data_out(8199) <= data_in(10036);
     data_out(8200) <= data_in(10037);
     data_out(8201) <= data_in(10041);
     data_out(8202) <= data_in(10044);
     data_out(8203) <= data_in(10045);
     data_out(8204) <= data_in(10048);
     data_out(8205) <= data_in(10050);
     data_out(8206) <= data_in(10055);
     data_out(8207) <= data_in(10056);
     data_out(8208) <= data_in(10057);
     data_out(8209) <= data_in(10058);
     data_out(8210) <= data_in(10059);
     data_out(8211) <= data_in(10063);
     data_out(8212) <= data_in(10067);
     data_out(8213) <= data_in(10069);
     data_out(8214) <= data_in(10071);
     data_out(8215) <= data_in(10076);
     data_out(8216) <= data_in(10077);
     data_out(8217) <= data_in(10082);
     data_out(8218) <= data_in(10085);
     data_out(8219) <= data_in(10090);
     data_out(8220) <= data_in(10097);
     data_out(8221) <= data_in(10099);
     data_out(8222) <= data_in(10100);
     data_out(8223) <= data_in(10101);
     data_out(8224) <= data_in(10105);
     data_out(8225) <= data_in(10107);
     data_out(8226) <= data_in(10109);
     data_out(8227) <= data_in(10110);
     data_out(8228) <= data_in(10111);
     data_out(8229) <= data_in(10114);
     data_out(8230) <= data_in(10117);
     data_out(8231) <= data_in(10121);
     data_out(8232) <= data_in(10124);
     data_out(8233) <= data_in(10125);
     data_out(8234) <= data_in(10127);
     data_out(8235) <= data_in(10128);
     data_out(8236) <= data_in(10133);
     data_out(8237) <= data_in(10134);
     data_out(8238) <= data_in(10135);
     data_out(8239) <= data_in(10136);
     data_out(8240) <= data_in(10146);
     data_out(8241) <= data_in(10147);
     data_out(8242) <= data_in(10148);
     data_out(8243) <= data_in(10149);
     data_out(8244) <= data_in(10150);
     data_out(8245) <= data_in(10154);
     data_out(8246) <= data_in(10155);
     data_out(8247) <= data_in(10156);
     data_out(8248) <= data_in(10157);
     data_out(8249) <= data_in(10159);
     data_out(8250) <= data_in(10160);
     data_out(8251) <= data_in(10161);
     data_out(8252) <= data_in(10162);
     data_out(8253) <= data_in(10163);
     data_out(8254) <= data_in(10166);
     data_out(8255) <= data_in(10167);
     data_out(8256) <= data_in(10168);
     data_out(8257) <= data_in(10169);
     data_out(8258) <= data_in(10170);
     data_out(8259) <= data_in(10174);
     data_out(8260) <= data_in(10175);
     data_out(8261) <= data_in(10176);
     data_out(8262) <= data_in(10178);
     data_out(8263) <= data_in(10183);
     data_out(8264) <= data_in(10184);
     data_out(8265) <= data_in(10185);
     data_out(8266) <= data_in(10190);
     data_out(8267) <= data_in(10191);
     data_out(8268) <= data_in(10192);
     data_out(8269) <= data_in(10193);
     data_out(8270) <= data_in(10195);
     data_out(8271) <= data_in(10196);
     data_out(8272) <= data_in(10197);
     data_out(8273) <= data_in(10201);
     data_out(8274) <= data_in(10202);
     data_out(8275) <= data_in(10211);
     data_out(8276) <= data_in(10212);
     data_out(8277) <= data_in(10213);
     data_out(8278) <= data_in(10215);
     data_out(8279) <= data_in(10217);
     data_out(8280) <= data_in(10221);
     data_out(8281) <= data_in(10226);
     data_out(8282) <= data_in(10233);
     data_out(8283) <= data_in(10236);
     data_out(8284) <= data_in(10237);
     data_out(8285) <= data_in(10238);
     data_out(8286) <= data_in(364);
     data_out(8287) <= data_in(441);
     data_out(8288) <= data_in(473);
     data_out(8289) <= data_in(600);
     data_out(8290) <= data_in(969);
     data_out(8291) <= data_in(1009);
     data_out(8292) <= data_in(1123);
     data_out(8293) <= data_in(1296);
     data_out(8294) <= data_in(1900);
     data_out(8295) <= data_in(2145);
     data_out(8296) <= data_in(2256);
     data_out(8297) <= data_in(2262);
     data_out(8298) <= data_in(2284);
     data_out(8299) <= data_in(2352);
     data_out(8300) <= data_in(2408);
     data_out(8301) <= data_in(2452);
     data_out(8302) <= data_in(2478);
     data_out(8303) <= data_in(2483);
     data_out(8304) <= data_in(2565);
     data_out(8305) <= data_in(2732);
     data_out(8306) <= data_in(2842);
     data_out(8307) <= data_in(2901);
     data_out(8308) <= data_in(3038);
     data_out(8309) <= data_in(3151);
     data_out(8310) <= data_in(3182);
     data_out(8311) <= data_in(3246);
     data_out(8312) <= data_in(3410);
     data_out(8313) <= data_in(3557);
     data_out(8314) <= data_in(3731);
     data_out(8315) <= data_in(3736);
     data_out(8316) <= data_in(3818);
     data_out(8317) <= data_in(4203);
     data_out(8318) <= data_in(4265);
     data_out(8319) <= data_in(4471);
     data_out(8320) <= data_in(4498);
     data_out(8321) <= data_in(4533);
     data_out(8322) <= data_in(4547);
     data_out(8323) <= data_in(4548);
     data_out(8324) <= data_in(4550);
     data_out(8325) <= data_in(4557);
     data_out(8326) <= data_in(4796);
     data_out(8327) <= data_in(4803);
     data_out(8328) <= data_in(4818);
     data_out(8329) <= data_in(4897);
     data_out(8330) <= data_in(4982);
     data_out(8331) <= data_in(4994);
     data_out(8332) <= data_in(5175);
     data_out(8333) <= data_in(5209);
     data_out(8334) <= data_in(5317);
     data_out(8335) <= data_in(6031);
     data_out(8336) <= data_in(6485);
     data_out(8337) <= data_in(6623);
     data_out(8338) <= data_in(6692);
     data_out(8339) <= data_in(7220);
     data_out(8340) <= data_in(7222);
     data_out(8341) <= data_in(7290);
     data_out(8342) <= data_in(7439);
     data_out(8343) <= data_in(7718);
     data_out(8344) <= data_in(8204);
     data_out(8345) <= data_in(8252);
     data_out(8346) <= data_in(8263);
     data_out(8347) <= data_in(8283);
     data_out(8348) <= data_in(8410);
     data_out(8349) <= data_in(8632);
     data_out(8350) <= data_in(8824);
     data_out(8351) <= data_in(8865);
     data_out(8352) <= data_in(8894);
     data_out(8353) <= data_in(9021);
     data_out(8354) <= data_in(9312);
     data_out(8355) <= data_in(9518);
     data_out(8356) <= data_in(9694);
     data_out(8357) <= data_in(9725);
     data_out(8358) <= data_in(9849);
     data_out(8359) <= data_in(9892);
     data_out(8360) <= data_in(10046);
     data_out(8361) <= data_in(10108);
     data_out(8362) <= data_in(562);
     data_out(8363) <= data_in(566);
     data_out(8364) <= data_in(669);
     data_out(8365) <= data_in(719);
     data_out(8366) <= data_in(1128);
     data_out(8367) <= data_in(1159);
     data_out(8368) <= data_in(1251);
     data_out(8369) <= data_in(1314);
     data_out(8370) <= data_in(1361);
     data_out(8371) <= data_in(1599);
     data_out(8372) <= data_in(1636);
     data_out(8373) <= data_in(1928);
     data_out(8374) <= data_in(2046);
     data_out(8375) <= data_in(2259);
     data_out(8376) <= data_in(2309);
     data_out(8377) <= data_in(2707);
     data_out(8378) <= data_in(2764);
     data_out(8379) <= data_in(2953);
     data_out(8380) <= data_in(2961);
     data_out(8381) <= data_in(3609);
     data_out(8382) <= data_in(3616);
     data_out(8383) <= data_in(3620);
     data_out(8384) <= data_in(4463);
     data_out(8385) <= data_in(4742);
     data_out(8386) <= data_in(4853);
     data_out(8387) <= data_in(5139);
     data_out(8388) <= data_in(5208);
     data_out(8389) <= data_in(5210);
     data_out(8390) <= data_in(5232);
     data_out(8391) <= data_in(5491);
     data_out(8392) <= data_in(6400);
     data_out(8393) <= data_in(6532);
     data_out(8394) <= data_in(6743);
     data_out(8395) <= data_in(6975);
     data_out(8396) <= data_in(7567);
     data_out(8397) <= data_in(7700);
     data_out(8398) <= data_in(7974);
     data_out(8399) <= data_in(8118);
     data_out(8400) <= data_in(8147);
     data_out(8401) <= data_in(8222);
     data_out(8402) <= data_in(8257);
     data_out(8403) <= data_in(8373);
     data_out(8404) <= data_in(8485);
     data_out(8405) <= data_in(8702);
     data_out(8406) <= data_in(8850);
     data_out(8407) <= data_in(9158);
     data_out(8408) <= data_in(9233);
     data_out(8409) <= data_in(9506);
     data_out(8410) <= data_in(9873);
     data_out(8411) <= data_in(9878);
     data_out(8412) <= data_in(960);
     data_out(8413) <= data_in(979);
     data_out(8414) <= data_in(1048);
     data_out(8415) <= data_in(1286);
     data_out(8416) <= data_in(1474);
     data_out(8417) <= data_in(1534);
     data_out(8418) <= data_in(1601);
     data_out(8419) <= data_in(1639);
     data_out(8420) <= data_in(1750);
     data_out(8421) <= data_in(1958);
     data_out(8422) <= data_in(2293);
     data_out(8423) <= data_in(2297);
     data_out(8424) <= data_in(2530);
     data_out(8425) <= data_in(2733);
     data_out(8426) <= data_in(2826);
     data_out(8427) <= data_in(2999);
     data_out(8428) <= data_in(3030);
     data_out(8429) <= data_in(3386);
     data_out(8430) <= data_in(3470);
     data_out(8431) <= data_in(3799);
     data_out(8432) <= data_in(4025);
     data_out(8433) <= data_in(4101);
     data_out(8434) <= data_in(4183);
     data_out(8435) <= data_in(4376);
     data_out(8436) <= data_in(4424);
     data_out(8437) <= data_in(4450);
     data_out(8438) <= data_in(4514);
     data_out(8439) <= data_in(4549);
     data_out(8440) <= data_in(4606);
     data_out(8441) <= data_in(4852);
     data_out(8442) <= data_in(4861);
     data_out(8443) <= data_in(4873);
     data_out(8444) <= data_in(5299);
     data_out(8445) <= data_in(5330);
     data_out(8446) <= data_in(5417);
     data_out(8447) <= data_in(5490);
     data_out(8448) <= data_in(5557);
     data_out(8449) <= data_in(5801);
     data_out(8450) <= data_in(6505);
     data_out(8451) <= data_in(6518);
     data_out(8452) <= data_in(6523);
     data_out(8453) <= data_in(6524);
     data_out(8454) <= data_in(6653);
     data_out(8455) <= data_in(6779);
     data_out(8456) <= data_in(6911);
     data_out(8457) <= data_in(6934);
     data_out(8458) <= data_in(7032);
     data_out(8459) <= data_in(7200);
     data_out(8460) <= data_in(7462);
     data_out(8461) <= data_in(7572);
     data_out(8462) <= data_in(7617);
     data_out(8463) <= data_in(7667);
     data_out(8464) <= data_in(7868);
     data_out(8465) <= data_in(7940);
     data_out(8466) <= data_in(8073);
     data_out(8467) <= data_in(8391);
     data_out(8468) <= data_in(8514);
     data_out(8469) <= data_in(8534);
     data_out(8470) <= data_in(8599);
     data_out(8471) <= data_in(8630);
     data_out(8472) <= data_in(8800);
     data_out(8473) <= data_in(9042);
     data_out(8474) <= data_in(9128);
     data_out(8475) <= data_in(9232);
     data_out(8476) <= data_in(9353);
     data_out(8477) <= data_in(9501);
     data_out(8478) <= data_in(9750);
     data_out(8479) <= data_in(9751);
     data_out(8480) <= data_in(10158);
     data_out(8481) <= data_in(10224);
     data_out(8482) <= data_in(424);
     data_out(8483) <= data_in(657);
     data_out(8484) <= data_in(764);
     data_out(8485) <= data_in(1042);
     data_out(8486) <= data_in(1375);
     data_out(8487) <= data_in(1462);
     data_out(8488) <= data_in(1465);
     data_out(8489) <= data_in(1505);
     data_out(8490) <= data_in(1934);
     data_out(8491) <= data_in(1993);
     data_out(8492) <= data_in(2425);
     data_out(8493) <= data_in(2501);
     data_out(8494) <= data_in(2690);
     data_out(8495) <= data_in(2759);
     data_out(8496) <= data_in(2785);
     data_out(8497) <= data_in(2985);
     data_out(8498) <= data_in(2994);
     data_out(8499) <= data_in(3146);
     data_out(8500) <= data_in(3245);
     data_out(8501) <= data_in(3333);
     data_out(8502) <= data_in(3356);
     data_out(8503) <= data_in(3520);
     data_out(8504) <= data_in(3614);
     data_out(8505) <= data_in(3726);
     data_out(8506) <= data_in(4018);
     data_out(8507) <= data_in(4170);
     data_out(8508) <= data_in(4209);
     data_out(8509) <= data_in(4347);
     data_out(8510) <= data_in(4355);
     data_out(8511) <= data_in(4365);
     data_out(8512) <= data_in(4604);
     data_out(8513) <= data_in(4634);
     data_out(8514) <= data_in(4648);
     data_out(8515) <= data_in(4834);
     data_out(8516) <= data_in(4886);
     data_out(8517) <= data_in(4960);
     data_out(8518) <= data_in(4980);
     data_out(8519) <= data_in(5016);
     data_out(8520) <= data_in(5073);
     data_out(8521) <= data_in(5095);
     data_out(8522) <= data_in(5101);
     data_out(8523) <= data_in(5189);
     data_out(8524) <= data_in(5307);
     data_out(8525) <= data_in(5366);
     data_out(8526) <= data_in(5612);
     data_out(8527) <= data_in(6231);
     data_out(8528) <= data_in(6236);
     data_out(8529) <= data_in(6345);
     data_out(8530) <= data_in(6662);
     data_out(8531) <= data_in(6792);
     data_out(8532) <= data_in(6904);
     data_out(8533) <= data_in(6992);
     data_out(8534) <= data_in(7008);
     data_out(8535) <= data_in(7194);
     data_out(8536) <= data_in(7234);
     data_out(8537) <= data_in(7419);
     data_out(8538) <= data_in(7716);
     data_out(8539) <= data_in(7754);
     data_out(8540) <= data_in(7811);
     data_out(8541) <= data_in(7944);
     data_out(8542) <= data_in(8119);
     data_out(8543) <= data_in(8154);
     data_out(8544) <= data_in(8206);
     data_out(8545) <= data_in(8423);
     data_out(8546) <= data_in(8503);
     data_out(8547) <= data_in(8882);
     data_out(8548) <= data_in(8935);
     data_out(8549) <= data_in(8983);
     data_out(8550) <= data_in(9073);
     data_out(8551) <= data_in(9270);
     data_out(8552) <= data_in(9359);
     data_out(8553) <= data_in(9389);
     data_out(8554) <= data_in(9418);
     data_out(8555) <= data_in(9823);
     data_out(8556) <= data_in(10033);
     data_out(8557) <= data_in(10227);
     data_out(8558) <= data_in(260);
     data_out(8559) <= data_in(261);
     data_out(8560) <= data_in(268);
     data_out(8561) <= data_in(283);
     data_out(8562) <= data_in(292);
     data_out(8563) <= data_in(417);
     data_out(8564) <= data_in(468);
     data_out(8565) <= data_in(483);
     data_out(8566) <= data_in(487);
     data_out(8567) <= data_in(567);
     data_out(8568) <= data_in(591);
     data_out(8569) <= data_in(732);
     data_out(8570) <= data_in(788);
     data_out(8571) <= data_in(830);
     data_out(8572) <= data_in(866);
     data_out(8573) <= data_in(916);
     data_out(8574) <= data_in(919);
     data_out(8575) <= data_in(931);
     data_out(8576) <= data_in(1031);
     data_out(8577) <= data_in(1093);
     data_out(8578) <= data_in(1105);
     data_out(8579) <= data_in(1169);
     data_out(8580) <= data_in(1240);
     data_out(8581) <= data_in(1244);
     data_out(8582) <= data_in(1331);
     data_out(8583) <= data_in(1392);
     data_out(8584) <= data_in(1402);
     data_out(8585) <= data_in(1430);
     data_out(8586) <= data_in(1451);
     data_out(8587) <= data_in(1461);
     data_out(8588) <= data_in(1488);
     data_out(8589) <= data_in(1494);
     data_out(8590) <= data_in(1588);
     data_out(8591) <= data_in(1757);
     data_out(8592) <= data_in(1810);
     data_out(8593) <= data_in(1813);
     data_out(8594) <= data_in(1884);
     data_out(8595) <= data_in(1935);
     data_out(8596) <= data_in(1970);
     data_out(8597) <= data_in(2005);
     data_out(8598) <= data_in(2011);
     data_out(8599) <= data_in(2059);
     data_out(8600) <= data_in(2124);
     data_out(8601) <= data_in(2164);
     data_out(8602) <= data_in(2176);
     data_out(8603) <= data_in(2223);
     data_out(8604) <= data_in(2253);
     data_out(8605) <= data_in(2320);
     data_out(8606) <= data_in(2347);
     data_out(8607) <= data_in(2376);
     data_out(8608) <= data_in(2377);
     data_out(8609) <= data_in(2417);
     data_out(8610) <= data_in(2442);
     data_out(8611) <= data_in(2528);
     data_out(8612) <= data_in(2586);
     data_out(8613) <= data_in(2610);
     data_out(8614) <= data_in(2618);
     data_out(8615) <= data_in(2662);
     data_out(8616) <= data_in(2944);
     data_out(8617) <= data_in(2957);
     data_out(8618) <= data_in(3039);
     data_out(8619) <= data_in(3084);
     data_out(8620) <= data_in(3160);
     data_out(8621) <= data_in(3177);
     data_out(8622) <= data_in(3236);
     data_out(8623) <= data_in(3242);
     data_out(8624) <= data_in(3379);
     data_out(8625) <= data_in(3569);
     data_out(8626) <= data_in(3673);
     data_out(8627) <= data_in(3709);
     data_out(8628) <= data_in(3873);
     data_out(8629) <= data_in(3901);
     data_out(8630) <= data_in(4002);
     data_out(8631) <= data_in(4016);
     data_out(8632) <= data_in(4197);
     data_out(8633) <= data_in(4268);
     data_out(8634) <= data_in(4290);
     data_out(8635) <= data_in(4313);
     data_out(8636) <= data_in(4320);
     data_out(8637) <= data_in(4322);
     data_out(8638) <= data_in(4328);
     data_out(8639) <= data_in(4366);
     data_out(8640) <= data_in(4390);
     data_out(8641) <= data_in(4431);
     data_out(8642) <= data_in(4488);
     data_out(8643) <= data_in(4563);
     data_out(8644) <= data_in(4787);
     data_out(8645) <= data_in(4821);
     data_out(8646) <= data_in(4830);
     data_out(8647) <= data_in(4839);
     data_out(8648) <= data_in(4926);
     data_out(8649) <= data_in(4981);
     data_out(8650) <= data_in(5055);
     data_out(8651) <= data_in(5086);
     data_out(8652) <= data_in(5213);
     data_out(8653) <= data_in(5238);
     data_out(8654) <= data_in(5379);
     data_out(8655) <= data_in(5422);
     data_out(8656) <= data_in(5450);
     data_out(8657) <= data_in(5468);
     data_out(8658) <= data_in(5480);
     data_out(8659) <= data_in(5493);
     data_out(8660) <= data_in(5601);
     data_out(8661) <= data_in(5622);
     data_out(8662) <= data_in(5679);
     data_out(8663) <= data_in(5686);
     data_out(8664) <= data_in(5709);
     data_out(8665) <= data_in(5844);
     data_out(8666) <= data_in(5860);
     data_out(8667) <= data_in(5899);
     data_out(8668) <= data_in(5935);
     data_out(8669) <= data_in(5973);
     data_out(8670) <= data_in(5988);
     data_out(8671) <= data_in(6044);
     data_out(8672) <= data_in(6048);
     data_out(8673) <= data_in(6054);
     data_out(8674) <= data_in(6102);
     data_out(8675) <= data_in(6117);
     data_out(8676) <= data_in(6167);
     data_out(8677) <= data_in(6235);
     data_out(8678) <= data_in(6295);
     data_out(8679) <= data_in(6598);
     data_out(8680) <= data_in(6611);
     data_out(8681) <= data_in(6614);
     data_out(8682) <= data_in(6729);
     data_out(8683) <= data_in(6769);
     data_out(8684) <= data_in(6790);
     data_out(8685) <= data_in(6822);
     data_out(8686) <= data_in(6836);
     data_out(8687) <= data_in(6873);
     data_out(8688) <= data_in(6956);
     data_out(8689) <= data_in(7102);
     data_out(8690) <= data_in(7109);
     data_out(8691) <= data_in(7120);
     data_out(8692) <= data_in(7148);
     data_out(8693) <= data_in(7244);
     data_out(8694) <= data_in(7264);
     data_out(8695) <= data_in(7303);
     data_out(8696) <= data_in(7310);
     data_out(8697) <= data_in(7314);
     data_out(8698) <= data_in(7359);
     data_out(8699) <= data_in(7422);
     data_out(8700) <= data_in(7444);
     data_out(8701) <= data_in(7478);
     data_out(8702) <= data_in(7512);
     data_out(8703) <= data_in(7558);
     data_out(8704) <= data_in(7560);
     data_out(8705) <= data_in(7620);
     data_out(8706) <= data_in(7633);
     data_out(8707) <= data_in(7639);
     data_out(8708) <= data_in(7683);
     data_out(8709) <= data_in(7710);
     data_out(8710) <= data_in(7711);
     data_out(8711) <= data_in(7752);
     data_out(8712) <= data_in(7834);
     data_out(8713) <= data_in(7920);
     data_out(8714) <= data_in(7933);
     data_out(8715) <= data_in(7936);
     data_out(8716) <= data_in(8113);
     data_out(8717) <= data_in(8198);
     data_out(8718) <= data_in(8231);
     data_out(8719) <= data_in(8234);
     data_out(8720) <= data_in(8238);
     data_out(8721) <= data_in(8287);
     data_out(8722) <= data_in(8324);
     data_out(8723) <= data_in(8365);
     data_out(8724) <= data_in(8396);
     data_out(8725) <= data_in(8461);
     data_out(8726) <= data_in(8561);
     data_out(8727) <= data_in(8619);
     data_out(8728) <= data_in(8637);
     data_out(8729) <= data_in(8821);
     data_out(8730) <= data_in(8863);
     data_out(8731) <= data_in(8984);
     data_out(8732) <= data_in(9025);
     data_out(8733) <= data_in(9083);
     data_out(8734) <= data_in(9137);
     data_out(8735) <= data_in(9191);
     data_out(8736) <= data_in(9211);
     data_out(8737) <= data_in(9214);
     data_out(8738) <= data_in(9243);
     data_out(8739) <= data_in(9390);
     data_out(8740) <= data_in(9442);
     data_out(8741) <= data_in(9588);
     data_out(8742) <= data_in(9794);
     data_out(8743) <= data_in(9856);
     data_out(8744) <= data_in(9865);
     data_out(8745) <= data_in(9877);
     data_out(8746) <= data_in(9969);
     data_out(8747) <= data_in(10015);
     data_out(8748) <= data_in(10034);
     data_out(8749) <= data_in(10064);
     data_out(8750) <= data_in(10116);
     data_out(8751) <= data_in(10189);
     data_out(8752) <= data_in(10208);
     data_out(8753) <= data_in(10222);
     data_out(8754) <= data_in(291);
     data_out(8755) <= data_in(524);
     data_out(8756) <= data_in(676);
     data_out(8757) <= data_in(895);
     data_out(8758) <= data_in(914);
     data_out(8759) <= data_in(975);
     data_out(8760) <= data_in(983);
     data_out(8761) <= data_in(1188);
     data_out(8762) <= data_in(1250);
     data_out(8763) <= data_in(1382);
     data_out(8764) <= data_in(1441);
     data_out(8765) <= data_in(1475);
     data_out(8766) <= data_in(1610);
     data_out(8767) <= data_in(1625);
     data_out(8768) <= data_in(1806);
     data_out(8769) <= data_in(1995);
     data_out(8770) <= data_in(2179);
     data_out(8771) <= data_in(2230);
     data_out(8772) <= data_in(2373);
     data_out(8773) <= data_in(2668);
     data_out(8774) <= data_in(2669);
     data_out(8775) <= data_in(2738);
     data_out(8776) <= data_in(2990);
     data_out(8777) <= data_in(3515);
     data_out(8778) <= data_in(3811);
     data_out(8779) <= data_in(3977);
     data_out(8780) <= data_in(4007);
     data_out(8781) <= data_in(4138);
     data_out(8782) <= data_in(4213);
     data_out(8783) <= data_in(4218);
     data_out(8784) <= data_in(4352);
     data_out(8785) <= data_in(4408);
     data_out(8786) <= data_in(4790);
     data_out(8787) <= data_in(4799);
     data_out(8788) <= data_in(4805);
     data_out(8789) <= data_in(5481);
     data_out(8790) <= data_in(5711);
     data_out(8791) <= data_in(5736);
     data_out(8792) <= data_in(5753);
     data_out(8793) <= data_in(6161);
     data_out(8794) <= data_in(6185);
     data_out(8795) <= data_in(6264);
     data_out(8796) <= data_in(6457);
     data_out(8797) <= data_in(6529);
     data_out(8798) <= data_in(6751);
     data_out(8799) <= data_in(6775);
     data_out(8800) <= data_in(7074);
     data_out(8801) <= data_in(7245);
     data_out(8802) <= data_in(7476);
     data_out(8803) <= data_in(7732);
     data_out(8804) <= data_in(7958);
     data_out(8805) <= data_in(8004);
     data_out(8806) <= data_in(8195);
     data_out(8807) <= data_in(8267);
     data_out(8808) <= data_in(8344);
     data_out(8809) <= data_in(8346);
     data_out(8810) <= data_in(8455);
     data_out(8811) <= data_in(8644);
     data_out(8812) <= data_in(9117);
     data_out(8813) <= data_in(9141);
     data_out(8814) <= data_in(9299);
     data_out(8815) <= data_in(9446);
     data_out(8816) <= data_in(9654);
     data_out(8817) <= data_in(9689);
     data_out(8818) <= data_in(10030);
     data_out(8819) <= data_in(10068);
     data_out(8820) <= data_in(10234);
     data_out(8821) <= data_in(249);
     data_out(8822) <= data_in(304);
     data_out(8823) <= data_in(319);
     data_out(8824) <= data_in(347);
     data_out(8825) <= data_in(387);
     data_out(8826) <= data_in(442);
     data_out(8827) <= data_in(445);
     data_out(8828) <= data_in(702);
     data_out(8829) <= data_in(706);
     data_out(8830) <= data_in(769);
     data_out(8831) <= data_in(862);
     data_out(8832) <= data_in(879);
     data_out(8833) <= data_in(893);
     data_out(8834) <= data_in(1013);
     data_out(8835) <= data_in(1110);
     data_out(8836) <= data_in(1158);
     data_out(8837) <= data_in(1226);
     data_out(8838) <= data_in(1295);
     data_out(8839) <= data_in(1297);
     data_out(8840) <= data_in(1352);
     data_out(8841) <= data_in(1444);
     data_out(8842) <= data_in(1492);
     data_out(8843) <= data_in(1542);
     data_out(8844) <= data_in(1562);
     data_out(8845) <= data_in(1565);
     data_out(8846) <= data_in(1658);
     data_out(8847) <= data_in(1710);
     data_out(8848) <= data_in(1774);
     data_out(8849) <= data_in(1826);
     data_out(8850) <= data_in(1835);
     data_out(8851) <= data_in(1864);
     data_out(8852) <= data_in(1921);
     data_out(8853) <= data_in(1952);
     data_out(8854) <= data_in(2008);
     data_out(8855) <= data_in(2096);
     data_out(8856) <= data_in(2097);
     data_out(8857) <= data_in(2172);
     data_out(8858) <= data_in(2193);
     data_out(8859) <= data_in(2304);
     data_out(8860) <= data_in(2378);
     data_out(8861) <= data_in(2381);
     data_out(8862) <= data_in(2428);
     data_out(8863) <= data_in(2486);
     data_out(8864) <= data_in(2489);
     data_out(8865) <= data_in(2500);
     data_out(8866) <= data_in(2545);
     data_out(8867) <= data_in(2567);
     data_out(8868) <= data_in(2652);
     data_out(8869) <= data_in(2656);
     data_out(8870) <= data_in(2689);
     data_out(8871) <= data_in(2693);
     data_out(8872) <= data_in(2702);
     data_out(8873) <= data_in(2749);
     data_out(8874) <= data_in(2767);
     data_out(8875) <= data_in(2894);
     data_out(8876) <= data_in(2918);
     data_out(8877) <= data_in(2929);
     data_out(8878) <= data_in(2977);
     data_out(8879) <= data_in(3025);
     data_out(8880) <= data_in(3169);
     data_out(8881) <= data_in(3189);
     data_out(8882) <= data_in(3305);
     data_out(8883) <= data_in(3312);
     data_out(8884) <= data_in(3347);
     data_out(8885) <= data_in(3364);
     data_out(8886) <= data_in(3373);
     data_out(8887) <= data_in(3404);
     data_out(8888) <= data_in(3544);
     data_out(8889) <= data_in(3593);
     data_out(8890) <= data_in(3641);
     data_out(8891) <= data_in(3757);
     data_out(8892) <= data_in(3760);
     data_out(8893) <= data_in(3774);
     data_out(8894) <= data_in(3777);
     data_out(8895) <= data_in(3813);
     data_out(8896) <= data_in(3890);
     data_out(8897) <= data_in(3926);
     data_out(8898) <= data_in(3937);
     data_out(8899) <= data_in(3988);
     data_out(8900) <= data_in(4060);
     data_out(8901) <= data_in(4062);
     data_out(8902) <= data_in(4085);
     data_out(8903) <= data_in(4149);
     data_out(8904) <= data_in(4150);
     data_out(8905) <= data_in(4169);
     data_out(8906) <= data_in(4172);
     data_out(8907) <= data_in(4194);
     data_out(8908) <= data_in(4281);
     data_out(8909) <= data_in(4486);
     data_out(8910) <= data_in(4493);
     data_out(8911) <= data_in(4502);
     data_out(8912) <= data_in(4506);
     data_out(8913) <= data_in(4544);
     data_out(8914) <= data_in(4572);
     data_out(8915) <= data_in(4593);
     data_out(8916) <= data_in(4603);
     data_out(8917) <= data_in(4743);
     data_out(8918) <= data_in(4786);
     data_out(8919) <= data_in(4850);
     data_out(8920) <= data_in(4884);
     data_out(8921) <= data_in(4935);
     data_out(8922) <= data_in(4971);
     data_out(8923) <= data_in(5193);
     data_out(8924) <= data_in(5202);
     data_out(8925) <= data_in(5410);
     data_out(8926) <= data_in(5465);
     data_out(8927) <= data_in(5485);
     data_out(8928) <= data_in(5664);
     data_out(8929) <= data_in(5723);
     data_out(8930) <= data_in(5768);
     data_out(8931) <= data_in(5786);
     data_out(8932) <= data_in(5806);
     data_out(8933) <= data_in(5807);
     data_out(8934) <= data_in(5983);
     data_out(8935) <= data_in(6017);
     data_out(8936) <= data_in(6164);
     data_out(8937) <= data_in(6166);
     data_out(8938) <= data_in(6220);
     data_out(8939) <= data_in(6246);
     data_out(8940) <= data_in(6307);
     data_out(8941) <= data_in(6460);
     data_out(8942) <= data_in(6555);
     data_out(8943) <= data_in(6561);
     data_out(8944) <= data_in(6602);
     data_out(8945) <= data_in(6698);
     data_out(8946) <= data_in(6723);
     data_out(8947) <= data_in(6732);
     data_out(8948) <= data_in(6889);
     data_out(8949) <= data_in(6915);
     data_out(8950) <= data_in(7028);
     data_out(8951) <= data_in(7031);
     data_out(8952) <= data_in(7040);
     data_out(8953) <= data_in(7096);
     data_out(8954) <= data_in(7205);
     data_out(8955) <= data_in(7227);
     data_out(8956) <= data_in(7316);
     data_out(8957) <= data_in(7369);
     data_out(8958) <= data_in(7423);
     data_out(8959) <= data_in(7498);
     data_out(8960) <= data_in(7540);
     data_out(8961) <= data_in(7600);
     data_out(8962) <= data_in(7610);
     data_out(8963) <= data_in(7638);
     data_out(8964) <= data_in(7736);
     data_out(8965) <= data_in(7829);
     data_out(8966) <= data_in(7873);
     data_out(8967) <= data_in(7891);
     data_out(8968) <= data_in(7895);
     data_out(8969) <= data_in(7899);
     data_out(8970) <= data_in(7904);
     data_out(8971) <= data_in(7932);
     data_out(8972) <= data_in(8001);
     data_out(8973) <= data_in(8013);
     data_out(8974) <= data_in(8191);
     data_out(8975) <= data_in(8200);
     data_out(8976) <= data_in(8219);
     data_out(8977) <= data_in(8228);
     data_out(8978) <= data_in(8266);
     data_out(8979) <= data_in(8308);
     data_out(8980) <= data_in(8478);
     data_out(8981) <= data_in(8578);
     data_out(8982) <= data_in(8715);
     data_out(8983) <= data_in(8757);
     data_out(8984) <= data_in(8985);
     data_out(8985) <= data_in(8999);
     data_out(8986) <= data_in(9024);
     data_out(8987) <= data_in(9032);
     data_out(8988) <= data_in(9091);
     data_out(8989) <= data_in(9177);
     data_out(8990) <= data_in(9241);
     data_out(8991) <= data_in(9300);
     data_out(8992) <= data_in(9342);
     data_out(8993) <= data_in(9454);
     data_out(8994) <= data_in(9476);
     data_out(8995) <= data_in(9559);
     data_out(8996) <= data_in(9573);
     data_out(8997) <= data_in(9596);
     data_out(8998) <= data_in(9612);
     data_out(8999) <= data_in(9671);
     data_out(9000) <= data_in(9726);
     data_out(9001) <= data_in(9733);
     data_out(9002) <= data_in(9793);
     data_out(9003) <= data_in(9826);
     data_out(9004) <= data_in(9830);
     data_out(9005) <= data_in(9896);
     data_out(9006) <= data_in(9922);
     data_out(9007) <= data_in(9934);
     data_out(9008) <= data_in(9994);
     data_out(9009) <= data_in(10143);
     data_out(9010) <= data_in(379);
     data_out(9011) <= data_in(609);
     data_out(9012) <= data_in(853);
     data_out(9013) <= data_in(932);
     data_out(9014) <= data_in(1269);
     data_out(9015) <= data_in(1379);
     data_out(9016) <= data_in(1403);
     data_out(9017) <= data_in(1535);
     data_out(9018) <= data_in(1815);
     data_out(9019) <= data_in(1965);
     data_out(9020) <= data_in(2485);
     data_out(9021) <= data_in(2513);
     data_out(9022) <= data_in(2722);
     data_out(9023) <= data_in(2742);
     data_out(9024) <= data_in(2962);
     data_out(9025) <= data_in(3268);
     data_out(9026) <= data_in(3406);
     data_out(9027) <= data_in(3463);
     data_out(9028) <= data_in(3524);
     data_out(9029) <= data_in(3531);
     data_out(9030) <= data_in(3552);
     data_out(9031) <= data_in(3788);
     data_out(9032) <= data_in(3970);
     data_out(9033) <= data_in(4109);
     data_out(9034) <= data_in(4199);
     data_out(9035) <= data_in(4325);
     data_out(9036) <= data_in(4387);
     data_out(9037) <= data_in(4527);
     data_out(9038) <= data_in(4591);
     data_out(9039) <= data_in(4841);
     data_out(9040) <= data_in(4965);
     data_out(9041) <= data_in(5587);
     data_out(9042) <= data_in(5989);
     data_out(9043) <= data_in(6091);
     data_out(9044) <= data_in(6153);
     data_out(9045) <= data_in(6271);
     data_out(9046) <= data_in(6386);
     data_out(9047) <= data_in(6462);
     data_out(9048) <= data_in(6789);
     data_out(9049) <= data_in(7100);
     data_out(9050) <= data_in(7146);
     data_out(9051) <= data_in(7158);
     data_out(9052) <= data_in(7283);
     data_out(9053) <= data_in(7388);
     data_out(9054) <= data_in(7534);
     data_out(9055) <= data_in(7569);
     data_out(9056) <= data_in(7570);
     data_out(9057) <= data_in(7580);
     data_out(9058) <= data_in(7801);
     data_out(9059) <= data_in(7844);
     data_out(9060) <= data_in(7896);
     data_out(9061) <= data_in(8092);
     data_out(9062) <= data_in(8165);
     data_out(9063) <= data_in(8321);
     data_out(9064) <= data_in(8372);
     data_out(9065) <= data_in(8940);
     data_out(9066) <= data_in(9015);
     data_out(9067) <= data_in(9075);
     data_out(9068) <= data_in(9311);
     data_out(9069) <= data_in(9498);
     data_out(9070) <= data_in(9504);
     data_out(9071) <= data_in(9507);
     data_out(9072) <= data_in(9532);
     data_out(9073) <= data_in(9715);
     data_out(9074) <= data_in(9757);
     data_out(9075) <= data_in(9779);
     data_out(9076) <= data_in(9796);
     data_out(9077) <= data_in(10001);
     data_out(9078) <= data_in(10087);
     data_out(9079) <= data_in(414);
     data_out(9080) <= data_in(444);
     data_out(9081) <= data_in(623);
     data_out(9082) <= data_in(870);
     data_out(9083) <= data_in(889);
     data_out(9084) <= data_in(994);
     data_out(9085) <= data_in(1162);
     data_out(9086) <= data_in(1293);
     data_out(9087) <= data_in(1307);
     data_out(9088) <= data_in(1691);
     data_out(9089) <= data_in(2119);
     data_out(9090) <= data_in(3059);
     data_out(9091) <= data_in(3123);
     data_out(9092) <= data_in(3323);
     data_out(9093) <= data_in(3415);
     data_out(9094) <= data_in(3729);
     data_out(9095) <= data_in(4587);
     data_out(9096) <= data_in(4683);
     data_out(9097) <= data_in(4707);
     data_out(9098) <= data_in(4813);
     data_out(9099) <= data_in(4997);
     data_out(9100) <= data_in(5142);
     data_out(9101) <= data_in(5224);
     data_out(9102) <= data_in(5405);
     data_out(9103) <= data_in(5473);
     data_out(9104) <= data_in(5577);
     data_out(9105) <= data_in(5617);
     data_out(9106) <= data_in(5696);
     data_out(9107) <= data_in(5726);
     data_out(9108) <= data_in(5747);
     data_out(9109) <= data_in(5832);
     data_out(9110) <= data_in(6150);
     data_out(9111) <= data_in(6412);
     data_out(9112) <= data_in(6442);
     data_out(9113) <= data_in(6563);
     data_out(9114) <= data_in(6685);
     data_out(9115) <= data_in(6741);
     data_out(9116) <= data_in(6839);
     data_out(9117) <= data_in(6886);
     data_out(9118) <= data_in(8101);
     data_out(9119) <= data_in(8157);
     data_out(9120) <= data_in(8174);
     data_out(9121) <= data_in(8311);
     data_out(9122) <= data_in(8378);
     data_out(9123) <= data_in(8399);
     data_out(9124) <= data_in(8405);
     data_out(9125) <= data_in(8494);
     data_out(9126) <= data_in(9003);
     data_out(9127) <= data_in(9009);
     data_out(9128) <= data_in(9189);
     data_out(9129) <= data_in(9296);
     data_out(9130) <= data_in(9426);
     data_out(9131) <= data_in(9468);
     data_out(9132) <= data_in(9481);
     data_out(9133) <= data_in(9541);
     data_out(9134) <= data_in(9548);
     data_out(9135) <= data_in(9621);
     data_out(9136) <= data_in(9837);
     data_out(9137) <= data_in(9859);
     data_out(9138) <= data_in(9868);
     data_out(9139) <= data_in(10179);
     data_out(9140) <= data_in(361);
     data_out(9141) <= data_in(1007);
     data_out(9142) <= data_in(1038);
     data_out(9143) <= data_in(1350);
     data_out(9144) <= data_in(1772);
     data_out(9145) <= data_in(1797);
     data_out(9146) <= data_in(1999);
     data_out(9147) <= data_in(2348);
     data_out(9148) <= data_in(2783);
     data_out(9149) <= data_in(2849);
     data_out(9150) <= data_in(3005);
     data_out(9151) <= data_in(3085);
     data_out(9152) <= data_in(3270);
     data_out(9153) <= data_in(3343);
     data_out(9154) <= data_in(3387);
     data_out(9155) <= data_in(3442);
     data_out(9156) <= data_in(3918);
     data_out(9157) <= data_in(4163);
     data_out(9158) <= data_in(4364);
     data_out(9159) <= data_in(4588);
     data_out(9160) <= data_in(4791);
     data_out(9161) <= data_in(4860);
     data_out(9162) <= data_in(5088);
     data_out(9163) <= data_in(5553);
     data_out(9164) <= data_in(5809);
     data_out(9165) <= data_in(6026);
     data_out(9166) <= data_in(6037);
     data_out(9167) <= data_in(6284);
     data_out(9168) <= data_in(6324);
     data_out(9169) <= data_in(6341);
     data_out(9170) <= data_in(6347);
     data_out(9171) <= data_in(6499);
     data_out(9172) <= data_in(6673);
     data_out(9173) <= data_in(6713);
     data_out(9174) <= data_in(6843);
     data_out(9175) <= data_in(6960);
     data_out(9176) <= data_in(6973);
     data_out(9177) <= data_in(7225);
     data_out(9178) <= data_in(7460);
     data_out(9179) <= data_in(7511);
     data_out(9180) <= data_in(7758);
     data_out(9181) <= data_in(8104);
     data_out(9182) <= data_in(8258);
     data_out(9183) <= data_in(8309);
     data_out(9184) <= data_in(8839);
     data_out(9185) <= data_in(8924);
     data_out(9186) <= data_in(9230);
     data_out(9187) <= data_in(9246);
     data_out(9188) <= data_in(9305);
     data_out(9189) <= data_in(9576);
     data_out(9190) <= data_in(295);
     data_out(9191) <= data_in(326);
     data_out(9192) <= data_in(502);
     data_out(9193) <= data_in(568);
     data_out(9194) <= data_in(678);
     data_out(9195) <= data_in(838);
     data_out(9196) <= data_in(1056);
     data_out(9197) <= data_in(1060);
     data_out(9198) <= data_in(1068);
     data_out(9199) <= data_in(1249);
     data_out(9200) <= data_in(1370);
     data_out(9201) <= data_in(1408);
     data_out(9202) <= data_in(1419);
     data_out(9203) <= data_in(1458);
     data_out(9204) <= data_in(1989);
     data_out(9205) <= data_in(2042);
     data_out(9206) <= data_in(3071);
     data_out(9207) <= data_in(3080);
     data_out(9208) <= data_in(3124);
     data_out(9209) <= data_in(3335);
     data_out(9210) <= data_in(3369);
     data_out(9211) <= data_in(3516);
     data_out(9212) <= data_in(3814);
     data_out(9213) <= data_in(3830);
     data_out(9214) <= data_in(4031);
     data_out(9215) <= data_in(4039);
     data_out(9216) <= data_in(4253);
     data_out(9217) <= data_in(4292);
     data_out(9218) <= data_in(4327);
     data_out(9219) <= data_in(4392);
     data_out(9220) <= data_in(4434);
     data_out(9221) <= data_in(4449);
     data_out(9222) <= data_in(5464);
     data_out(9223) <= data_in(5749);
     data_out(9224) <= data_in(5755);
     data_out(9225) <= data_in(5850);
     data_out(9226) <= data_in(5885);
     data_out(9227) <= data_in(6130);
     data_out(9228) <= data_in(6309);
     data_out(9229) <= data_in(6469);
     data_out(9230) <= data_in(6484);
     data_out(9231) <= data_in(6500);
     data_out(9232) <= data_in(6872);
     data_out(9233) <= data_in(6946);
     data_out(9234) <= data_in(6953);
     data_out(9235) <= data_in(6970);
     data_out(9236) <= data_in(7179);
     data_out(9237) <= data_in(7259);
     data_out(9238) <= data_in(7272);
     data_out(9239) <= data_in(7308);
     data_out(9240) <= data_in(7712);
     data_out(9241) <= data_in(7846);
     data_out(9242) <= data_in(8025);
     data_out(9243) <= data_in(8034);
     data_out(9244) <= data_in(8259);
     data_out(9245) <= data_in(8339);
     data_out(9246) <= data_in(8362);
     data_out(9247) <= data_in(8635);
     data_out(9248) <= data_in(8646);
     data_out(9249) <= data_in(8667);
     data_out(9250) <= data_in(8756);
     data_out(9251) <= data_in(8786);
     data_out(9252) <= data_in(9430);
     data_out(9253) <= data_in(9525);
     data_out(9254) <= data_in(9939);
     data_out(9255) <= data_in(257);
     data_out(9256) <= data_in(362);
     data_out(9257) <= data_in(372);
     data_out(9258) <= data_in(556);
     data_out(9259) <= data_in(923);
     data_out(9260) <= data_in(946);
     data_out(9261) <= data_in(1126);
     data_out(9262) <= data_in(1256);
     data_out(9263) <= data_in(1261);
     data_out(9264) <= data_in(1274);
     data_out(9265) <= data_in(1291);
     data_out(9266) <= data_in(1907);
     data_out(9267) <= data_in(1985);
     data_out(9268) <= data_in(2072);
     data_out(9269) <= data_in(2226);
     data_out(9270) <= data_in(2701);
     data_out(9271) <= data_in(2839);
     data_out(9272) <= data_in(2896);
     data_out(9273) <= data_in(2963);
     data_out(9274) <= data_in(3092);
     data_out(9275) <= data_in(3199);
     data_out(9276) <= data_in(3546);
     data_out(9277) <= data_in(3745);
     data_out(9278) <= data_in(4076);
     data_out(9279) <= data_in(4093);
     data_out(9280) <= data_in(4748);
     data_out(9281) <= data_in(5132);
     data_out(9282) <= data_in(5173);
     data_out(9283) <= data_in(5456);
     data_out(9284) <= data_in(5602);
     data_out(9285) <= data_in(5910);
     data_out(9286) <= data_in(6055);
     data_out(9287) <= data_in(6109);
     data_out(9288) <= data_in(6325);
     data_out(9289) <= data_in(6463);
     data_out(9290) <= data_in(6553);
     data_out(9291) <= data_in(6749);
     data_out(9292) <= data_in(6996);
     data_out(9293) <= data_in(7045);
     data_out(9294) <= data_in(7630);
     data_out(9295) <= data_in(7848);
     data_out(9296) <= data_in(7987);
     data_out(9297) <= data_in(8058);
     data_out(9298) <= data_in(8242);
     data_out(9299) <= data_in(8395);
     data_out(9300) <= data_in(8448);
     data_out(9301) <= data_in(8507);
     data_out(9302) <= data_in(8620);
     data_out(9303) <= data_in(8673);
     data_out(9304) <= data_in(8742);
     data_out(9305) <= data_in(8867);
     data_out(9306) <= data_in(8973);
     data_out(9307) <= data_in(9245);
     data_out(9308) <= data_in(9308);
     data_out(9309) <= data_in(9396);
     data_out(9310) <= data_in(9408);
     data_out(9311) <= data_in(9916);
     data_out(9312) <= data_in(10054);
     data_out(9313) <= data_in(290);
     data_out(9314) <= data_in(320);
     data_out(9315) <= data_in(493);
     data_out(9316) <= data_in(639);
     data_out(9317) <= data_in(736);
     data_out(9318) <= data_in(737);
     data_out(9319) <= data_in(997);
     data_out(9320) <= data_in(1163);
     data_out(9321) <= data_in(1294);
     data_out(9322) <= data_in(1341);
     data_out(9323) <= data_in(1418);
     data_out(9324) <= data_in(1843);
     data_out(9325) <= data_in(1918);
     data_out(9326) <= data_in(2128);
     data_out(9327) <= data_in(2225);
     data_out(9328) <= data_in(2308);
     data_out(9329) <= data_in(2334);
     data_out(9330) <= data_in(2337);
     data_out(9331) <= data_in(2644);
     data_out(9332) <= data_in(2645);
     data_out(9333) <= data_in(2773);
     data_out(9334) <= data_in(2791);
     data_out(9335) <= data_in(2823);
     data_out(9336) <= data_in(3032);
     data_out(9337) <= data_in(3176);
     data_out(9338) <= data_in(3252);
     data_out(9339) <= data_in(3340);
     data_out(9340) <= data_in(3604);
     data_out(9341) <= data_in(3605);
     data_out(9342) <= data_in(3655);
     data_out(9343) <= data_in(3949);
     data_out(9344) <= data_in(4034);
     data_out(9345) <= data_in(4175);
     data_out(9346) <= data_in(4326);
     data_out(9347) <= data_in(4671);
     data_out(9348) <= data_in(4679);
     data_out(9349) <= data_in(4717);
     data_out(9350) <= data_in(4929);
     data_out(9351) <= data_in(5156);
     data_out(9352) <= data_in(5225);
     data_out(9353) <= data_in(5397);
     data_out(9354) <= data_in(5424);
     data_out(9355) <= data_in(5440);
     data_out(9356) <= data_in(5623);
     data_out(9357) <= data_in(5647);
     data_out(9358) <= data_in(5656);
     data_out(9359) <= data_in(5790);
     data_out(9360) <= data_in(5793);
     data_out(9361) <= data_in(5919);
     data_out(9362) <= data_in(5964);
     data_out(9363) <= data_in(5966);
     data_out(9364) <= data_in(5984);
     data_out(9365) <= data_in(6021);
     data_out(9366) <= data_in(6063);
     data_out(9367) <= data_in(6100);
     data_out(9368) <= data_in(6108);
     data_out(9369) <= data_in(6186);
     data_out(9370) <= data_in(6230);
     data_out(9371) <= data_in(6430);
     data_out(9372) <= data_in(6450);
     data_out(9373) <= data_in(6691);
     data_out(9374) <= data_in(6813);
     data_out(9375) <= data_in(7073);
     data_out(9376) <= data_in(7301);
     data_out(9377) <= data_in(7463);
     data_out(9378) <= data_in(7516);
     data_out(9379) <= data_in(7526);
     data_out(9380) <= data_in(7657);
     data_out(9381) <= data_in(7786);
     data_out(9382) <= data_in(7905);
     data_out(9383) <= data_in(7976);
     data_out(9384) <= data_in(8094);
     data_out(9385) <= data_in(8235);
     data_out(9386) <= data_in(8488);
     data_out(9387) <= data_in(8708);
     data_out(9388) <= data_in(8990);
     data_out(9389) <= data_in(9065);
     data_out(9390) <= data_in(9144);
     data_out(9391) <= data_in(9159);
     data_out(9392) <= data_in(9491);
     data_out(9393) <= data_in(9539);
     data_out(9394) <= data_in(9584);
     data_out(9395) <= data_in(9840);
     data_out(9396) <= data_in(9853);
     data_out(9397) <= data_in(9951);
     data_out(9398) <= data_in(9954);
     data_out(9399) <= data_in(10006);
     data_out(9400) <= data_in(10016);
     data_out(9401) <= data_in(10089);
     data_out(9402) <= data_in(10140);
     data_out(9403) <= data_in(10194);
     data_out(9404) <= data_in(10231);
     data_out(9405) <= data_in(620);
     data_out(9406) <= data_in(1028);
     data_out(9407) <= data_in(1311);
     data_out(9408) <= data_in(1329);
     data_out(9409) <= data_in(1496);
     data_out(9410) <= data_in(1852);
     data_out(9411) <= data_in(1877);
     data_out(9412) <= data_in(2057);
     data_out(9413) <= data_in(2058);
     data_out(9414) <= data_in(2149);
     data_out(9415) <= data_in(2370);
     data_out(9416) <= data_in(2579);
     data_out(9417) <= data_in(2598);
     data_out(9418) <= data_in(2741);
     data_out(9419) <= data_in(2857);
     data_out(9420) <= data_in(3075);
     data_out(9421) <= data_in(3353);
     data_out(9422) <= data_in(3389);
     data_out(9423) <= data_in(3566);
     data_out(9424) <= data_in(3972);
     data_out(9425) <= data_in(4491);
     data_out(9426) <= data_in(4908);
     data_out(9427) <= data_in(4936);
     data_out(9428) <= data_in(5573);
     data_out(9429) <= data_in(5965);
     data_out(9430) <= data_in(6042);
     data_out(9431) <= data_in(6112);
     data_out(9432) <= data_in(6320);
     data_out(9433) <= data_in(6331);
     data_out(9434) <= data_in(6366);
     data_out(9435) <= data_in(6865);
     data_out(9436) <= data_in(7018);
     data_out(9437) <= data_in(7024);
     data_out(9438) <= data_in(7086);
     data_out(9439) <= data_in(7161);
     data_out(9440) <= data_in(7250);
     data_out(9441) <= data_in(7344);
     data_out(9442) <= data_in(7433);
     data_out(9443) <= data_in(7650);
     data_out(9444) <= data_in(7750);
     data_out(9445) <= data_in(7912);
     data_out(9446) <= data_in(7950);
     data_out(9447) <= data_in(8591);
     data_out(9448) <= data_in(8594);
     data_out(9449) <= data_in(8945);
     data_out(9450) <= data_in(8993);
     data_out(9451) <= data_in(9652);
     data_out(9452) <= data_in(9702);
     data_out(9453) <= data_in(10129);
     data_out(9454) <= data_in(10223);
     data_out(9455) <= data_in(271);
     data_out(9456) <= data_in(331);
     data_out(9457) <= data_in(391);
     data_out(9458) <= data_in(535);
     data_out(9459) <= data_in(748);
     data_out(9460) <= data_in(781);
     data_out(9461) <= data_in(815);
     data_out(9462) <= data_in(841);
     data_out(9463) <= data_in(910);
     data_out(9464) <= data_in(913);
     data_out(9465) <= data_in(936);
     data_out(9466) <= data_in(940);
     data_out(9467) <= data_in(963);
     data_out(9468) <= data_in(972);
     data_out(9469) <= data_in(1087);
     data_out(9470) <= data_in(1320);
     data_out(9471) <= data_in(1482);
     data_out(9472) <= data_in(1580);
     data_out(9473) <= data_in(1817);
     data_out(9474) <= data_in(1941);
     data_out(9475) <= data_in(2024);
     data_out(9476) <= data_in(2114);
     data_out(9477) <= data_in(2416);
     data_out(9478) <= data_in(2445);
     data_out(9479) <= data_in(2801);
     data_out(9480) <= data_in(3094);
     data_out(9481) <= data_in(3319);
     data_out(9482) <= data_in(3334);
     data_out(9483) <= data_in(3416);
     data_out(9484) <= data_in(3485);
     data_out(9485) <= data_in(3602);
     data_out(9486) <= data_in(3762);
     data_out(9487) <= data_in(3771);
     data_out(9488) <= data_in(3787);
     data_out(9489) <= data_in(3807);
     data_out(9490) <= data_in(3944);
     data_out(9491) <= data_in(3947);
     data_out(9492) <= data_in(3997);
     data_out(9493) <= data_in(4023);
     data_out(9494) <= data_in(4053);
     data_out(9495) <= data_in(4058);
     data_out(9496) <= data_in(4153);
     data_out(9497) <= data_in(4189);
     data_out(9498) <= data_in(4407);
     data_out(9499) <= data_in(4627);
     data_out(9500) <= data_in(4642);
     data_out(9501) <= data_in(4670);
     data_out(9502) <= data_in(4833);
     data_out(9503) <= data_in(4851);
     data_out(9504) <= data_in(5153);
     data_out(9505) <= data_in(5212);
     data_out(9506) <= data_in(5296);
     data_out(9507) <= data_in(5743);
     data_out(9508) <= data_in(5909);
     data_out(9509) <= data_in(6086);
     data_out(9510) <= data_in(6209);
     data_out(9511) <= data_in(6380);
     data_out(9512) <= data_in(6719);
     data_out(9513) <= data_in(6851);
     data_out(9514) <= data_in(7112);
     data_out(9515) <= data_in(7135);
     data_out(9516) <= data_in(7180);
     data_out(9517) <= data_in(7186);
     data_out(9518) <= data_in(7187);
     data_out(9519) <= data_in(7281);
     data_out(9520) <= data_in(7405);
     data_out(9521) <= data_in(7581);
     data_out(9522) <= data_in(7818);
     data_out(9523) <= data_in(8074);
     data_out(9524) <= data_in(8098);
     data_out(9525) <= data_in(8145);
     data_out(9526) <= data_in(8812);
     data_out(9527) <= data_in(8969);
     data_out(9528) <= data_in(8998);
     data_out(9529) <= data_in(9074);
     data_out(9530) <= data_in(9115);
     data_out(9531) <= data_in(9179);
     data_out(9532) <= data_in(9229);
     data_out(9533) <= data_in(9264);
     data_out(9534) <= data_in(9301);
     data_out(9535) <= data_in(9326);
     data_out(9536) <= data_in(9329);
     data_out(9537) <= data_in(9457);
     data_out(9538) <= data_in(9574);
     data_out(9539) <= data_in(9643);
     data_out(9540) <= data_in(9744);
     data_out(9541) <= data_in(9924);
     data_out(9542) <= data_in(9977);
     data_out(9543) <= data_in(10123);
     data_out(9544) <= data_in(10239);
     data_out(9545) <= data_in(447);
     data_out(9546) <= data_in(452);
     data_out(9547) <= data_in(671);
     data_out(9548) <= data_in(1062);
     data_out(9549) <= data_in(1145);
     data_out(9550) <= data_in(1543);
     data_out(9551) <= data_in(1577);
     data_out(9552) <= data_in(1994);
     data_out(9553) <= data_in(2103);
     data_out(9554) <= data_in(2178);
     data_out(9555) <= data_in(2307);
     data_out(9556) <= data_in(2628);
     data_out(9557) <= data_in(2725);
     data_out(9558) <= data_in(2888);
     data_out(9559) <= data_in(3083);
     data_out(9560) <= data_in(3223);
     data_out(9561) <= data_in(3226);
     data_out(9562) <= data_in(3509);
     data_out(9563) <= data_in(3556);
     data_out(9564) <= data_in(3963);
     data_out(9565) <= data_in(3992);
     data_out(9566) <= data_in(4121);
     data_out(9567) <= data_in(4357);
     data_out(9568) <= data_in(4462);
     data_out(9569) <= data_in(4831);
     data_out(9570) <= data_in(5454);
     data_out(9571) <= data_in(5996);
     data_out(9572) <= data_in(6299);
     data_out(9573) <= data_in(6403);
     data_out(9574) <= data_in(7053);
     data_out(9575) <= data_in(7645);
     data_out(9576) <= data_in(7663);
     data_out(9577) <= data_in(7858);
     data_out(9578) <= data_in(8122);
     data_out(9579) <= data_in(8273);
     data_out(9580) <= data_in(8282);
     data_out(9581) <= data_in(8294);
     data_out(9582) <= data_in(8490);
     data_out(9583) <= data_in(8556);
     data_out(9584) <= data_in(8895);
     data_out(9585) <= data_in(8965);
     data_out(9586) <= data_in(9317);
     data_out(9587) <= data_in(9394);
     data_out(9588) <= data_in(9527);
     data_out(9589) <= data_in(9831);
     data_out(9590) <= data_in(9836);
     data_out(9591) <= data_in(10043);
     data_out(9592) <= data_in(286);
     data_out(9593) <= data_in(881);
     data_out(9594) <= data_in(1040);
     data_out(9595) <= data_in(1052);
     data_out(9596) <= data_in(1164);
     data_out(9597) <= data_in(1196);
     data_out(9598) <= data_in(1455);
     data_out(9599) <= data_in(1516);
     data_out(9600) <= data_in(1803);
     data_out(9601) <= data_in(1976);
     data_out(9602) <= data_in(2167);
     data_out(9603) <= data_in(2245);
     data_out(9604) <= data_in(2584);
     data_out(9605) <= data_in(2633);
     data_out(9606) <= data_in(2697);
     data_out(9607) <= data_in(2915);
     data_out(9608) <= data_in(2968);
     data_out(9609) <= data_in(3004);
     data_out(9610) <= data_in(3103);
     data_out(9611) <= data_in(3363);
     data_out(9612) <= data_in(3527);
     data_out(9613) <= data_in(3668);
     data_out(9614) <= data_in(3698);
     data_out(9615) <= data_in(3816);
     data_out(9616) <= data_in(3826);
     data_out(9617) <= data_in(3916);
     data_out(9618) <= data_in(3925);
     data_out(9619) <= data_in(4009);
     data_out(9620) <= data_in(4090);
     data_out(9621) <= data_in(4104);
     data_out(9622) <= data_in(4239);
     data_out(9623) <= data_in(4577);
     data_out(9624) <= data_in(4721);
     data_out(9625) <= data_in(5058);
     data_out(9626) <= data_in(5161);
     data_out(9627) <= data_in(5275);
     data_out(9628) <= data_in(5294);
     data_out(9629) <= data_in(5302);
     data_out(9630) <= data_in(5371);
     data_out(9631) <= data_in(5517);
     data_out(9632) <= data_in(5645);
     data_out(9633) <= data_in(5902);
     data_out(9634) <= data_in(6315);
     data_out(9635) <= data_in(6510);
     data_out(9636) <= data_in(6527);
     data_out(9637) <= data_in(6588);
     data_out(9638) <= data_in(6777);
     data_out(9639) <= data_in(6965);
     data_out(9640) <= data_in(7182);
     data_out(9641) <= data_in(7198);
     data_out(9642) <= data_in(7389);
     data_out(9643) <= data_in(7865);
     data_out(9644) <= data_in(7923);
     data_out(9645) <= data_in(7931);
     data_out(9646) <= data_in(8138);
     data_out(9647) <= data_in(8616);
     data_out(9648) <= data_in(8905);
     data_out(9649) <= data_in(9008);
     data_out(9650) <= data_in(9226);
     data_out(9651) <= data_in(9332);
     data_out(9652) <= data_in(9378);
     data_out(9653) <= data_in(9395);
     data_out(9654) <= data_in(9443);
     data_out(9655) <= data_in(9625);
     data_out(9656) <= data_in(9678);
     data_out(9657) <= data_in(9775);
     data_out(9658) <= data_in(9910);
     data_out(9659) <= data_in(9946);
     data_out(9660) <= data_in(9997);
     data_out(9661) <= data_in(10088);
     data_out(9662) <= data_in(334);
     data_out(9663) <= data_in(428);
     data_out(9664) <= data_in(602);
     data_out(9665) <= data_in(613);
     data_out(9666) <= data_in(1023);
     data_out(9667) <= data_in(1281);
     data_out(9668) <= data_in(1409);
     data_out(9669) <= data_in(1416);
     data_out(9670) <= data_in(1429);
     data_out(9671) <= data_in(1574);
     data_out(9672) <= data_in(1607);
     data_out(9673) <= data_in(1784);
     data_out(9674) <= data_in(1825);
     data_out(9675) <= data_in(2204);
     data_out(9676) <= data_in(2254);
     data_out(9677) <= data_in(2336);
     data_out(9678) <= data_in(2423);
     data_out(9679) <= data_in(2476);
     data_out(9680) <= data_in(2692);
     data_out(9681) <= data_in(2789);
     data_out(9682) <= data_in(3064);
     data_out(9683) <= data_in(3143);
     data_out(9684) <= data_in(3325);
     data_out(9685) <= data_in(3424);
     data_out(9686) <= data_in(3462);
     data_out(9687) <= data_in(3503);
     data_out(9688) <= data_in(3675);
     data_out(9689) <= data_in(3885);
     data_out(9690) <= data_in(4084);
     data_out(9691) <= data_in(4214);
     data_out(9692) <= data_in(4280);
     data_out(9693) <= data_in(4307);
     data_out(9694) <= data_in(4874);
     data_out(9695) <= data_in(5077);
     data_out(9696) <= data_in(5162);
     data_out(9697) <= data_in(5310);
     data_out(9698) <= data_in(5499);
     data_out(9699) <= data_in(5663);
     data_out(9700) <= data_in(5802);
     data_out(9701) <= data_in(6201);
     data_out(9702) <= data_in(6716);
     data_out(9703) <= data_in(6914);
     data_out(9704) <= data_in(7107);
     data_out(9705) <= data_in(7601);
     data_out(9706) <= data_in(7734);
     data_out(9707) <= data_in(7794);
     data_out(9708) <= data_in(7914);
     data_out(9709) <= data_in(7915);
     data_out(9710) <= data_in(8298);
     data_out(9711) <= data_in(8359);
     data_out(9712) <= data_in(8445);
     data_out(9713) <= data_in(8463);
     data_out(9714) <= data_in(8483);
     data_out(9715) <= data_in(8508);
     data_out(9716) <= data_in(8545);
     data_out(9717) <= data_in(8577);
     data_out(9718) <= data_in(8709);
     data_out(9719) <= data_in(8927);
     data_out(9720) <= data_in(9112);
     data_out(9721) <= data_in(9380);
     data_out(9722) <= data_in(9472);
     data_out(9723) <= data_in(9493);
     data_out(9724) <= data_in(9515);
     data_out(9725) <= data_in(9614);
     data_out(9726) <= data_in(9639);
     data_out(9727) <= data_in(9699);
     data_out(9728) <= data_in(9844);
     data_out(9729) <= data_in(9894);
     data_out(9730) <= data_in(9907);
     data_out(9731) <= data_in(311);
     data_out(9732) <= data_in(322);
     data_out(9733) <= data_in(349);
     data_out(9734) <= data_in(593);
     data_out(9735) <= data_in(677);
     data_out(9736) <= data_in(744);
     data_out(9737) <= data_in(773);
     data_out(9738) <= data_in(837);
     data_out(9739) <= data_in(938);
     data_out(9740) <= data_in(961);
     data_out(9741) <= data_in(1047);
     data_out(9742) <= data_in(1053);
     data_out(9743) <= data_in(1058);
     data_out(9744) <= data_in(1113);
     data_out(9745) <= data_in(1114);
     data_out(9746) <= data_in(1197);
     data_out(9747) <= data_in(1317);
     data_out(9748) <= data_in(1359);
     data_out(9749) <= data_in(1395);
     data_out(9750) <= data_in(1423);
     data_out(9751) <= data_in(1446);
     data_out(9752) <= data_in(1526);
     data_out(9753) <= data_in(1550);
     data_out(9754) <= data_in(1554);
     data_out(9755) <= data_in(1579);
     data_out(9756) <= data_in(1647);
     data_out(9757) <= data_in(1655);
     data_out(9758) <= data_in(1931);
     data_out(9759) <= data_in(1936);
     data_out(9760) <= data_in(2044);
     data_out(9761) <= data_in(2111);
     data_out(9762) <= data_in(2211);
     data_out(9763) <= data_in(2346);
     data_out(9764) <= data_in(2435);
     data_out(9765) <= data_in(2469);
     data_out(9766) <= data_in(2554);
     data_out(9767) <= data_in(2557);
     data_out(9768) <= data_in(2619);
     data_out(9769) <= data_in(2623);
     data_out(9770) <= data_in(2700);
     data_out(9771) <= data_in(2723);
     data_out(9772) <= data_in(2833);
     data_out(9773) <= data_in(2854);
     data_out(9774) <= data_in(2949);
     data_out(9775) <= data_in(3119);
     data_out(9776) <= data_in(3141);
     data_out(9777) <= data_in(3285);
     data_out(9778) <= data_in(3654);
     data_out(9779) <= data_in(3693);
     data_out(9780) <= data_in(3705);
     data_out(9781) <= data_in(3938);
     data_out(9782) <= data_in(3987);
     data_out(9783) <= data_in(4041);
     data_out(9784) <= data_in(4045);
     data_out(9785) <= data_in(4066);
     data_out(9786) <= data_in(4206);
     data_out(9787) <= data_in(4367);
     data_out(9788) <= data_in(4444);
     data_out(9789) <= data_in(4611);
     data_out(9790) <= data_in(4669);
     data_out(9791) <= data_in(4766);
     data_out(9792) <= data_in(4989);
     data_out(9793) <= data_in(4998);
     data_out(9794) <= data_in(5017);
     data_out(9795) <= data_in(5127);
     data_out(9796) <= data_in(5129);
     data_out(9797) <= data_in(5200);
     data_out(9798) <= data_in(5352);
     data_out(9799) <= data_in(5412);
     data_out(9800) <= data_in(5467);
     data_out(9801) <= data_in(5492);
     data_out(9802) <= data_in(5767);
     data_out(9803) <= data_in(5769);
     data_out(9804) <= data_in(5800);
     data_out(9805) <= data_in(5810);
     data_out(9806) <= data_in(5849);
     data_out(9807) <= data_in(5933);
     data_out(9808) <= data_in(6045);
     data_out(9809) <= data_in(6061);
     data_out(9810) <= data_in(6092);
     data_out(9811) <= data_in(6096);
     data_out(9812) <= data_in(6154);
     data_out(9813) <= data_in(6158);
     data_out(9814) <= data_in(6162);
     data_out(9815) <= data_in(6348);
     data_out(9816) <= data_in(6350);
     data_out(9817) <= data_in(6387);
     data_out(9818) <= data_in(6515);
     data_out(9819) <= data_in(6517);
     data_out(9820) <= data_in(6810);
     data_out(9821) <= data_in(6875);
     data_out(9822) <= data_in(6918);
     data_out(9823) <= data_in(6944);
     data_out(9824) <= data_in(7094);
     data_out(9825) <= data_in(7155);
     data_out(9826) <= data_in(7176);
     data_out(9827) <= data_in(7251);
     data_out(9828) <= data_in(7438);
     data_out(9829) <= data_in(7491);
     data_out(9830) <= data_in(7783);
     data_out(9831) <= data_in(7795);
     data_out(9832) <= data_in(7941);
     data_out(9833) <= data_in(8009);
     data_out(9834) <= data_in(8063);
     data_out(9835) <= data_in(8146);
     data_out(9836) <= data_in(8207);
     data_out(9837) <= data_in(8360);
     data_out(9838) <= data_in(8464);
     data_out(9839) <= data_in(8526);
     data_out(9840) <= data_in(8568);
     data_out(9841) <= data_in(8586);
     data_out(9842) <= data_in(8738);
     data_out(9843) <= data_in(8740);
     data_out(9844) <= data_in(8771);
     data_out(9845) <= data_in(8775);
     data_out(9846) <= data_in(8936);
     data_out(9847) <= data_in(8956);
     data_out(9848) <= data_in(9051);
     data_out(9849) <= data_in(9093);
     data_out(9850) <= data_in(9420);
     data_out(9851) <= data_in(9447);
     data_out(9852) <= data_in(9645);
     data_out(9853) <= data_in(9687);
     data_out(9854) <= data_in(10137);
     data_out(9855) <= data_in(10144);
     data_out(9856) <= data_in(282);
     data_out(9857) <= data_in(594);
     data_out(9858) <= data_in(603);
     data_out(9859) <= data_in(755);
     data_out(9860) <= data_in(1177);
     data_out(9861) <= data_in(1189);
     data_out(9862) <= data_in(1337);
     data_out(9863) <= data_in(1481);
     data_out(9864) <= data_in(1811);
     data_out(9865) <= data_in(1967);
     data_out(9866) <= data_in(1968);
     data_out(9867) <= data_in(1977);
     data_out(9868) <= data_in(2107);
     data_out(9869) <= data_in(2232);
     data_out(9870) <= data_in(2345);
     data_out(9871) <= data_in(2664);
     data_out(9872) <= data_in(2667);
     data_out(9873) <= data_in(3104);
     data_out(9874) <= data_in(3194);
     data_out(9875) <= data_in(3302);
     data_out(9876) <= data_in(3310);
     data_out(9877) <= data_in(3450);
     data_out(9878) <= data_in(3915);
     data_out(9879) <= data_in(3928);
     data_out(9880) <= data_in(4052);
     data_out(9881) <= data_in(4343);
     data_out(9882) <= data_in(4428);
     data_out(9883) <= data_in(4451);
     data_out(9884) <= data_in(4552);
     data_out(9885) <= data_in(4629);
     data_out(9886) <= data_in(4730);
     data_out(9887) <= data_in(4806);
     data_out(9888) <= data_in(4815);
     data_out(9889) <= data_in(4951);
     data_out(9890) <= data_in(4992);
     data_out(9891) <= data_in(5026);
     data_out(9892) <= data_in(5044);
     data_out(9893) <= data_in(5215);
     data_out(9894) <= data_in(5391);
     data_out(9895) <= data_in(5961);
     data_out(9896) <= data_in(6127);
     data_out(9897) <= data_in(6244);
     data_out(9898) <= data_in(6526);
     data_out(9899) <= data_in(6567);
     data_out(9900) <= data_in(6923);
     data_out(9901) <= data_in(7027);
     data_out(9902) <= data_in(7276);
     data_out(9903) <= data_in(7503);
     data_out(9904) <= data_in(7685);
     data_out(9905) <= data_in(7747);
     data_out(9906) <= data_in(7888);
     data_out(9907) <= data_in(7954);
     data_out(9908) <= data_in(8652);
     data_out(9909) <= data_in(8674);
     data_out(9910) <= data_in(8760);
     data_out(9911) <= data_in(8902);
     data_out(9912) <= data_in(8912);
     data_out(9913) <= data_in(9027);
     data_out(9914) <= data_in(9071);
     data_out(9915) <= data_in(9200);
     data_out(9916) <= data_in(9399);
     data_out(9917) <= data_in(9656);
     data_out(9918) <= data_in(9846);
     data_out(9919) <= data_in(9903);
     data_out(9920) <= data_in(9928);
     data_out(9921) <= data_in(9948);
     data_out(9922) <= data_in(9978);
     data_out(9923) <= data_in(243);
     data_out(9924) <= data_in(528);
     data_out(9925) <= data_in(534);
     data_out(9926) <= data_in(776);
     data_out(9927) <= data_in(1021);
     data_out(9928) <= data_in(1615);
     data_out(9929) <= data_in(2194);
     data_out(9930) <= data_in(2471);
     data_out(9931) <= data_in(2940);
     data_out(9932) <= data_in(3653);
     data_out(9933) <= data_in(4621);
     data_out(9934) <= data_in(5021);
     data_out(9935) <= data_in(5121);
     data_out(9936) <= data_in(5483);
     data_out(9937) <= data_in(5539);
     data_out(9938) <= data_in(5636);
     data_out(9939) <= data_in(5924);
     data_out(9940) <= data_in(6015);
     data_out(9941) <= data_in(6292);
     data_out(9942) <= data_in(6571);
     data_out(9943) <= data_in(6683);
     data_out(9944) <= data_in(6858);
     data_out(9945) <= data_in(7051);
     data_out(9946) <= data_in(7221);
     data_out(9947) <= data_in(7312);
     data_out(9948) <= data_in(7656);
     data_out(9949) <= data_in(8230);
     data_out(9950) <= data_in(8511);
     data_out(9951) <= data_in(8553);
     data_out(9952) <= data_in(8722);
     data_out(9953) <= data_in(8744);
     data_out(9954) <= data_in(8966);
     data_out(9955) <= data_in(9023);
     data_out(9956) <= data_in(9777);
     data_out(9957) <= data_in(9956);
     data_out(9958) <= data_in(10005);
     data_out(9959) <= data_in(10092);
     data_out(9960) <= data_in(10232);
     data_out(9961) <= data_in(356);
     data_out(9962) <= data_in(437);
     data_out(9963) <= data_in(541);
     data_out(9964) <= data_in(656);
     data_out(9965) <= data_in(1078);
     data_out(9966) <= data_in(1094);
     data_out(9967) <= data_in(1181);
     data_out(9968) <= data_in(1330);
     data_out(9969) <= data_in(1438);
     data_out(9970) <= data_in(1522);
     data_out(9971) <= data_in(1807);
     data_out(9972) <= data_in(1829);
     data_out(9973) <= data_in(1950);
     data_out(9974) <= data_in(2069);
     data_out(9975) <= data_in(2491);
     data_out(9976) <= data_in(2592);
     data_out(9977) <= data_in(2710);
     data_out(9978) <= data_in(2739);
     data_out(9979) <= data_in(3135);
     data_out(9980) <= data_in(3301);
     data_out(9981) <= data_in(3441);
     data_out(9982) <= data_in(3792);
     data_out(9983) <= data_in(3820);
     data_out(9984) <= data_in(4132);
     data_out(9985) <= data_in(4266);
     data_out(9986) <= data_in(4592);
     data_out(9987) <= data_in(4848);
     data_out(9988) <= data_in(4912);
     data_out(9989) <= data_in(5186);
     data_out(9990) <= data_in(5351);
     data_out(9991) <= data_in(5523);
     data_out(9992) <= data_in(5624);
     data_out(9993) <= data_in(5694);
     data_out(9994) <= data_in(5922);
     data_out(9995) <= data_in(5929);
     data_out(9996) <= data_in(6071);
     data_out(9997) <= data_in(6124);
     data_out(9998) <= data_in(6453);
     data_out(9999) <= data_in(6584);
     data_out(10000) <= data_in(6612);
     data_out(10001) <= data_in(6841);
     data_out(10002) <= data_in(7269);
     data_out(10003) <= data_in(7406);
     data_out(10004) <= data_in(7676);
     data_out(10005) <= data_in(7773);
     data_out(10006) <= data_in(7799);
     data_out(10007) <= data_in(8091);
     data_out(10008) <= data_in(8190);
     data_out(10009) <= data_in(8486);
     data_out(10010) <= data_in(8651);
     data_out(10011) <= data_in(8729);
     data_out(10012) <= data_in(8897);
     data_out(10013) <= data_in(8900);
     data_out(10014) <= data_in(8947);
     data_out(10015) <= data_in(9172);
     data_out(10016) <= data_in(9344);
     data_out(10017) <= data_in(9444);
     data_out(10018) <= data_in(9471);
     data_out(10019) <= data_in(9477);
     data_out(10020) <= data_in(9522);
     data_out(10021) <= data_in(9538);
     data_out(10022) <= data_in(9597);
     data_out(10023) <= data_in(9633);
     data_out(10024) <= data_in(9665);
     data_out(10025) <= data_in(9669);
     data_out(10026) <= data_in(9763);
     data_out(10027) <= data_in(9778);
     data_out(10028) <= data_in(9995);
     data_out(10029) <= data_in(783);
     data_out(10030) <= data_in(1050);
     data_out(10031) <= data_in(1530);
     data_out(10032) <= data_in(1714);
     data_out(10033) <= data_in(1910);
     data_out(10034) <= data_in(2197);
     data_out(10035) <= data_in(2339);
     data_out(10036) <= data_in(2821);
     data_out(10037) <= data_in(3263);
     data_out(10038) <= data_in(3506);
     data_out(10039) <= data_in(3583);
     data_out(10040) <= data_in(3878);
     data_out(10041) <= data_in(3982);
     data_out(10042) <= data_in(4382);
     data_out(10043) <= data_in(4404);
     data_out(10044) <= data_in(4802);
     data_out(10045) <= data_in(4876);
     data_out(10046) <= data_in(5134);
     data_out(10047) <= data_in(5306);
     data_out(10048) <= data_in(5355);
     data_out(10049) <= data_in(5678);
     data_out(10050) <= data_in(5861);
     data_out(10051) <= data_in(5963);
     data_out(10052) <= data_in(6099);
     data_out(10053) <= data_in(6379);
     data_out(10054) <= data_in(7077);
     data_out(10055) <= data_in(7121);
     data_out(10056) <= data_in(7211);
     data_out(10057) <= data_in(7223);
     data_out(10058) <= data_in(7692);
     data_out(10059) <= data_in(8418);
     data_out(10060) <= data_in(8475);
     data_out(10061) <= data_in(8567);
     data_out(10062) <= data_in(8779);
     data_out(10063) <= data_in(8830);
     data_out(10064) <= data_in(8877);
     data_out(10065) <= data_in(9040);
     data_out(10066) <= data_in(9708);
     data_out(10067) <= data_in(10130);
     data_out(10068) <= data_in(10220);
     data_out(10069) <= data_in(480);
     data_out(10070) <= data_in(514);
     data_out(10071) <= data_in(630);
     data_out(10072) <= data_in(642);
     data_out(10073) <= data_in(683);
     data_out(10074) <= data_in(791);
     data_out(10075) <= data_in(1010);
     data_out(10076) <= data_in(1241);
     data_out(10077) <= data_in(1514);
     data_out(10078) <= data_in(1740);
     data_out(10079) <= data_in(2227);
     data_out(10080) <= data_in(2450);
     data_out(10081) <= data_in(2480);
     data_out(10082) <= data_in(2712);
     data_out(10083) <= data_in(2730);
     data_out(10084) <= data_in(2864);
     data_out(10085) <= data_in(3196);
     data_out(10086) <= data_in(3464);
     data_out(10087) <= data_in(3730);
     data_out(10088) <= data_in(4143);
     data_out(10089) <= data_in(4151);
     data_out(10090) <= data_in(4160);
     data_out(10091) <= data_in(4258);
     data_out(10092) <= data_in(4701);
     data_out(10093) <= data_in(4855);
     data_out(10094) <= data_in(5039);
     data_out(10095) <= data_in(5148);
     data_out(10096) <= data_in(5194);
     data_out(10097) <= data_in(5507);
     data_out(10098) <= data_in(5575);
     data_out(10099) <= data_in(5611);
     data_out(10100) <= data_in(5764);
     data_out(10101) <= data_in(6179);
     data_out(10102) <= data_in(6558);
     data_out(10103) <= data_in(6835);
     data_out(10104) <= data_in(7149);
     data_out(10105) <= data_in(7203);
     data_out(10106) <= data_in(7260);
     data_out(10107) <= data_in(7317);
     data_out(10108) <= data_in(7383);
     data_out(10109) <= data_in(7494);
     data_out(10110) <= data_in(7603);
     data_out(10111) <= data_in(7708);
     data_out(10112) <= data_in(7751);
     data_out(10113) <= data_in(7837);
     data_out(10114) <= data_in(7911);
     data_out(10115) <= data_in(8015);
     data_out(10116) <= data_in(8057);
     data_out(10117) <= data_in(8107);
     data_out(10118) <= data_in(8213);
     data_out(10119) <= data_in(8442);
     data_out(10120) <= data_in(8558);
     data_out(10121) <= data_in(8719);
     data_out(10122) <= data_in(8762);
     data_out(10123) <= data_in(8881);
     data_out(10124) <= data_in(9068);
     data_out(10125) <= data_in(9404);
     data_out(10126) <= data_in(9598);
     data_out(10127) <= data_in(9670);
     data_out(10128) <= data_in(9747);
     data_out(10129) <= data_in(9827);
     data_out(10130) <= data_in(9984);
     data_out(10131) <= data_in(10024);
     data_out(10132) <= data_in(280);
     data_out(10133) <= data_in(314);
     data_out(10134) <= data_in(378);
     data_out(10135) <= data_in(771);
     data_out(10136) <= data_in(806);
     data_out(10137) <= data_in(810);
     data_out(10138) <= data_in(823);
     data_out(10139) <= data_in(848);
     data_out(10140) <= data_in(1018);
     data_out(10141) <= data_in(1143);
     data_out(10142) <= data_in(1316);
     data_out(10143) <= data_in(1343);
     data_out(10144) <= data_in(1490);
     data_out(10145) <= data_in(1544);
     data_out(10146) <= data_in(1559);
     data_out(10147) <= data_in(1560);
     data_out(10148) <= data_in(1597);
     data_out(10149) <= data_in(1649);
     data_out(10150) <= data_in(1889);
     data_out(10151) <= data_in(1981);
     data_out(10152) <= data_in(2115);
     data_out(10153) <= data_in(2594);
     data_out(10154) <= data_in(2673);
     data_out(10155) <= data_in(2792);
     data_out(10156) <= data_in(2934);
     data_out(10157) <= data_in(3018);
     data_out(10158) <= data_in(3026);
     data_out(10159) <= data_in(3029);
     data_out(10160) <= data_in(3035);
     data_out(10161) <= data_in(3042);
     data_out(10162) <= data_in(3049);
     data_out(10163) <= data_in(3057);
     data_out(10164) <= data_in(3063);
     data_out(10165) <= data_in(3109);
     data_out(10166) <= data_in(3167);
     data_out(10167) <= data_in(3296);
     data_out(10168) <= data_in(3390);
     data_out(10169) <= data_in(3486);
     data_out(10170) <= data_in(3577);
     data_out(10171) <= data_in(3893);
     data_out(10172) <= data_in(3995);
     data_out(10173) <= data_in(4050);
     data_out(10174) <= data_in(4222);
     data_out(10175) <= data_in(4238);
     data_out(10176) <= data_in(4248);
     data_out(10177) <= data_in(4262);
     data_out(10178) <= data_in(4291);
     data_out(10179) <= data_in(4323);
     data_out(10180) <= data_in(4371);
     data_out(10181) <= data_in(4525);
     data_out(10182) <= data_in(4555);
     data_out(10183) <= data_in(4673);
     data_out(10184) <= data_in(4749);
     data_out(10185) <= data_in(4811);
     data_out(10186) <= data_in(4974);
     data_out(10187) <= data_in(5009);
     data_out(10188) <= data_in(5203);
     data_out(10189) <= data_in(5222);
     data_out(10190) <= data_in(5266);
     data_out(10191) <= data_in(5335);
     data_out(10192) <= data_in(5358);
     data_out(10193) <= data_in(5364);
     data_out(10194) <= data_in(5515);
     data_out(10195) <= data_in(5737);
     data_out(10196) <= data_in(5745);
     data_out(10197) <= data_in(5782);
     data_out(10198) <= data_in(5866);
     data_out(10199) <= data_in(6303);
     data_out(10200) <= data_in(6312);
     data_out(10201) <= data_in(6432);
     data_out(10202) <= data_in(6445);
     data_out(10203) <= data_in(6474);
     data_out(10204) <= data_in(6599);
     data_out(10205) <= data_in(6639);
     data_out(10206) <= data_in(6781);
     data_out(10207) <= data_in(6796);
     data_out(10208) <= data_in(6831);
     data_out(10209) <= data_in(6912);
     data_out(10210) <= data_in(6930);
     data_out(10211) <= data_in(6931);
     data_out(10212) <= data_in(7029);
     data_out(10213) <= data_in(7527);
     data_out(10214) <= data_in(7660);
     data_out(10215) <= data_in(7702);
     data_out(10216) <= data_in(7797);
     data_out(10217) <= data_in(7831);
     data_out(10218) <= data_in(8186);
     data_out(10219) <= data_in(8436);
     data_out(10220) <= data_in(8438);
     data_out(10221) <= data_in(8454);
     data_out(10222) <= data_in(8467);
     data_out(10223) <= data_in(8498);
     data_out(10224) <= data_in(8736);
     data_out(10225) <= data_in(8752);
     data_out(10226) <= data_in(8778);
     data_out(10227) <= data_in(8845);
     data_out(10228) <= data_in(8861);
     data_out(10229) <= data_in(9111);
     data_out(10230) <= data_in(9171);
     data_out(10231) <= data_in(9248);
     data_out(10232) <= data_in(9540);
     data_out(10233) <= data_in(9629);
     data_out(10234) <= data_in(9674);
     data_out(10235) <= data_in(9790);
     data_out(10236) <= data_in(9807);
     data_out(10237) <= data_in(9891);
     data_out(10238) <= data_in(9933);
     data_out(10239) <= data_in(10091);
end Behavioral;



----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


entity reading_counter is
    generic (
        dimension_size     : integer := 1024;   -- dimension size 
        dimension_WIDTH    : integer := 10;     -- log2 dimension size 
        class_size    : integer := 10;     -- number of classes
        ECC_WIDTH          : integer := 8       -- bit-width of ECC_code 
    );
	port (
	clk                     : in std_logic;
    rst                     : in std_logic;
	din 					: in std_logic_vector(dimension_size-1 downto 0);
    count_reg               : in std_logic_vector(dimension_WIDTH-1 downto 0);
    dout                    : out std_logic_vector(dimension_WIDTH-1 downto 0)
	);	
end entity;

architecture behavior of reading_counter is

    -- Array types
    type CHV_memory_array is array (0 to dimension_size-1) of std_logic_vector(class_size-1 downto 0);
    type countingCheck is array (0 to dimension_WIDTH-1) of std_logic_vector(dimension_WIDTH-1 downto 0);

    -- Signals
    signal CHV_memory               : CHV_memory_array;
    signal CHV_memory_out : std_logic_vector(class_size-1 downto 0);
    signal corrected_CHV_memory_out : std_logic_vector(class_size-1 downto 0);
	signal din_suffle 					: std_logic_vector(dimension_size-1 downto 0);

    signal count_sim               : countingCheck;
    signal double_error    : std_logic;

    -- File I/O
    
    signal en_pops_regular         : std_logic_vector(class_size-1 downto 0);
    
    signal LFSRasHVCheck           : std_logic;
    signal LFSR_suffleAsHVCheck    : std_logic;

	signal ECC_out             : std_logic_vector(5-1 downto 0);
    
begin

    CHVMem: entity work.CHV_mem_10000
    port map(
        clk  => clk,
        address => count_reg,
        data => CHV_memory_out
    );

    HVmapper: entity work.dic_mapper 
    generic map(WIDTH => dimension_size)
    port map(
        data_in => din,
        data_out => din_suffle
    );

	ECCuut: entity work.ECC_vhdl_module
    generic map(
        C  => class_size,
        ECC_bit => 5   )
    port map(
        d => CHV_memory_out,
        p => ECC_out,
        double_error => double_error,
        dcw   => corrected_CHV_memory_out
    );
    
	ECCuutMem: entity work.configurable_counter
    generic map(
        dimension_WIDTH    =>  dimension_WIDTH,
        ECC_WIDTH => ECC_WIDTH   )
    port map(
        clk  => clk,
        rst  => rst,
        CHV_pointer => count_reg,
        ECC_out => ECC_out
    );

    LFSRasHVCheck  <= din_suffle(to_integer(unsigned(count_reg)));

    en_regular_pops: for k in 0 to class_size-1 generate
        en_pops_regular(k) <= corrected_CHV_memory_out(k) xor LFSRasHVCheck;
    end generate;

    -- Counters for regular
    class_counter: for k in 0 to class_size-1 generate
        simcounter: entity work.popCount 
            generic map(lenPop => dimension_WIDTH)
            port map(
                clk  => clk,
                rst  => rst,
                en   => en_pops_regular(k),
                dout => count_sim(k)
            );
    end generate;
	
	dout <= std_logic_vector(unsigned(count_sim(0)) + unsigned(count_sim(1)) + unsigned(count_sim(2)) + unsigned(count_sim(3)) + unsigned(count_sim(4)) + unsigned(count_sim(5)) + unsigned(count_sim(6)) + unsigned(count_sim(7)) + unsigned(count_sim(8)) + unsigned(count_sim(9)));
end architecture;



