

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ECC_vhdl_module is
    generic (
        C      : integer := 10;        -- Bit width number of classes or the segments size that we are going to correct
        ECC_bit: integer := 5          -- Number of bits for correction each column
    );
    port (
        d           : in  std_logic_vector(C-1 downto 0);  -- Input data vector
        p           : in  std_logic_vector(ECC_bit-1 downto 0);  -- Input ECC bits
        double_error: out std_logic;                        -- Output flag for double error
        dcw         : out std_logic_vector(C-1 downto 0)    -- Corrected data vector
    );
	attribute DONT_TOUCH : string;
	attribute KEEP : string;
	attribute DONT_TOUCH of ECC_vhdl_module : entity is "TRUE";
	attribute KEEP of ECC_vhdl_module : entity is "TRUE";
end entity ECC_vhdl_module;

architecture Behavioral of ECC_vhdl_module is
    signal dp : std_logic_vector(4 downto 0);  -- Parity calculated from input data
    signal s  : std_logic_vector(4 downto 0);  -- Syndrome bits
    signal df : std_logic_vector(9 downto 0);  -- Flag bit for getting correct data
    signal xw : std_logic;                     -- Intermediate signal for double error flag
begin

    -- Data Parity calculation
    dp(0) <= d(0) xor d(1) xor d(3) xor d(4) xor d(6) xor d(8);
    dp(1) <= d(0) xor d(2) xor d(3) xor d(5) xor d(6) xor d(9);
    dp(2) <= d(1) xor d(2) xor d(3) xor d(7) xor d(8) xor d(9);
    dp(3) <= d(4) xor d(5) xor d(6) xor d(7) xor d(8) xor d(9);
    dp(4) <= d(0) xor d(1) xor d(2) xor d(3) xor d(4) xor d(5) xor d(6) xor d(7) xor d(8) xor d(9) xor p(0) xor p(1) xor p(2) xor p(3);

    -- Syndrome: xor with actual parity
    s(0) <= p(0) xor dp(0);
    s(1) <= p(1) xor dp(1);
    s(2) <= p(2) xor dp(2);
    s(3) <= p(3) xor dp(3);
    s(4) <= p(4) xor dp(4);

    -- Flag bit for getting correct data
    df(0) <= s(0) and s(1) and not s(2) and not s(3) and s(4);
    df(1) <= s(0) and not s(1) and s(2) and not s(3) and s(4);
    df(2) <= not s(0) and s(1) and s(2) and not s(3) and s(4);
    df(3) <= s(0) and s(1) and s(2) and not s(3) and s(4);
    df(4) <= s(0) and not s(1) and not s(2) and s(3) and s(4);
    df(5) <= not s(0) and s(1) and not s(2) and s(3) and s(4);
    df(6) <= s(0) and s(1) and not s(2) and s(3) and s(4);
    df(7) <= not s(0) and not s(1) and s(2) and s(3) and s(4);
    df(8) <= s(0) and not s(1) and s(2) and s(3) and s(4);
    df(9) <= not s(0) and s(1) and s(2) and s(3) and s(4);

    -- Corrected data bits
    dcw(0) <= df(0) xor d(0);
    dcw(1) <= df(1) xor d(1);
    dcw(2) <= df(2) xor d(2);
    dcw(3) <= df(3) xor d(3);
    dcw(4) <= df(4) xor d(4);
    dcw(5) <= df(5) xor d(5);
    dcw(6) <= df(6) xor d(6);
    dcw(7) <= df(7) xor d(7);
    dcw(8) <= df(8) xor d(8);
    dcw(9) <= df(9) xor d(9);

    -- Intermediate signal for double error flag
    xw <= s(0) or s(1) or s(2) or s(3);

    -- Flag for double error
    double_error <= not s(4) and xw;  -- If 1, that means double error exists

end architecture Behavioral;


---------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY popCount IS
	GENERIC (lenPop : INTEGER := 8);   -- bit width out popCounters --- LOG2(#feature)
	PORT (
		clk , rst 	: IN STD_LOGIC;
		en		 	: IN STD_LOGIC;
		dout        : OUT  STD_LOGIC_VECTOR (lenPop-1 DOWNTO 0)
	);
	attribute DONT_TOUCH : string;
	attribute KEEP : string;
	attribute DONT_TOUCH of popCount : entity is "TRUE";
	attribute KEEP of popCount : entity is "TRUE";
END ENTITY popCount;

ARCHITECTURE behavioral OF popCount IS
SIGNAL popOut : STD_LOGIC_VECTOR (lenPop - 1 DOWNTO 0);
	
BEGIN

	PROCESS(clk)
		BEGIN 
		    IF rising_edge(clk) THEN
			    IF(rst = '1')THEN
				   popOut <= (OTHERS=>'0');
				ELSIF (en ='1') THEN 
				   popOut <= STD_LOGIC_VECTOR (UNSIGNED(popOut) + 1);
				END IF;
			END IF;
	END PROCESS;

	dout <= popOut;
END ARCHITECTURE behavioral;

---------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CHV_mem_10000 is
    Port (
        clk     : in  STD_LOGIC;
        address : in  STD_LOGIC_VECTOR(13 downto 0);
        data    : out STD_LOGIC_VECTOR(10 downto 0)
    );
end CHV_mem_10000;

architecture Behavioral of CHV_mem_10000 is
begin
    process(clk)
    begin
        if rising_edge(clk) then
            case address is
                when x"00" => data <= "1010110001";
                when x"01" => data <= "0100000000";
                when x"02" => data <= "0010101000";
                when x"03" => data <= "0100000000";
                when x"04" => data <= "1001010000";
                when x"05" => data <= "1011011011";
                when x"06" => data <= "0100000000";
                when x"07" => data <= "0100000000";
                when x"08" => data <= "0100000000";
                when x"09" => data <= "0010101000";
                when x"0A" => data <= "1110100111";
                when x"0B" => data <= "0100000000";
                when x"0C" => data <= "0100000000";
                when x"0D" => data <= "1001010000";
                when x"0E" => data <= "0100000000";
                when x"0F" => data <= "0100000000";
                when x"10" => data <= "0100110101";
                when x"11" => data <= "1111111000";
                when x"12" => data <= "1001010000";
                when x"13" => data <= "0100000000";
                when x"14" => data <= "1010000100";
                when x"15" => data <= "1011011011";
                when x"16" => data <= "0100000000";
                when x"17" => data <= "0100000000";
                when x"18" => data <= "0100000000";
                when x"19" => data <= "0100000000";
                when x"1A" => data <= "0100000000";
                when x"1B" => data <= "0011000010";
                when x"1C" => data <= "0100000000";
                when x"1D" => data <= "1001010000";
                when x"1E" => data <= "0100000000";
                when x"1F" => data <= "1000111010";
                when x"20" => data <= "0100000000";
                when x"21" => data <= "0100000000";
                when x"22" => data <= "0000100011";
                when x"23" => data <= "0100000000";
                when x"24" => data <= "0100000000";
                when x"25" => data <= "0100000000";
                when x"26" => data <= "1001010000";
                when x"27" => data <= "0100000000";
                when x"28" => data <= "0100000000";
                when x"29" => data <= "0100000000";
                when x"2A" => data <= "0100000000";
                when x"2B" => data <= "0100000000";
                when x"2C" => data <= "1001010000";
                when x"2D" => data <= "0100110101";
                when x"2E" => data <= "0100000000";
                when x"2F" => data <= "0100000000";
                when x"30" => data <= "0100000000";
                when x"31" => data <= "0100000000";
                when x"32" => data <= "0011000010";
                when x"33" => data <= "0100000000";
                when x"34" => data <= "0100000000";
                when x"35" => data <= "1001010000";
                when x"36" => data <= "0100000000";
                when x"37" => data <= "1001010000";
                when x"38" => data <= "0101011111";
                when x"39" => data <= "1001010000";
                when x"3A" => data <= "0100000000";
                when x"3B" => data <= "0110001011";
                when x"3C" => data <= "0100000000";
                when x"3D" => data <= "1110010010";
                when x"3E" => data <= "0100000000";
                when x"3F" => data <= "0101011111";
                when x"40" => data <= "0100000000";
                when x"41" => data <= "1010000100";
                when x"42" => data <= "0100000000";
                when x"43" => data <= "1111001101";
                when x"44" => data <= "0100000000";
                when x"45" => data <= "0100000000";
                when x"46" => data <= "0100000000";
                when x"47" => data <= "0100000000";
                when x"48" => data <= "0100110101";
                when x"49" => data <= "0100000000";
                when x"4A" => data <= "0011000010";
                when x"4B" => data <= "0100000000";
                when x"4C" => data <= "0100000000";
                when x"4D" => data <= "0100000000";
                when x"4E" => data <= "1101000110";
                when x"4F" => data <= "0100000000";
                when x"50" => data <= "1001010000";
                when x"51" => data <= "0100110101";
                when x"52" => data <= "0100000000";
                when x"53" => data <= "0100000000";
                when x"54" => data <= "0111100001";
                when x"55" => data <= "0100000000";
                when x"56" => data <= "1001010000";
                when x"57" => data <= "0100000000";
                when x"58" => data <= "0100000000";
                when x"59" => data <= "1110100111";
                when x"5A" => data <= "0100000000";
                when x"5B" => data <= "0010101000";
                when x"5C" => data <= "0100000000";
                when x"5D" => data <= "0100000000";
                when x"5E" => data <= "0100110101";
                when x"5F" => data <= "0100110101";
                when x"60" => data <= "0100000000";
                when x"61" => data <= "0100000000";
                when x"62" => data <= "0100000000";
                when x"63" => data <= "0100000000";
                when x"64" => data <= "1111111000";
                when x"65" => data <= "0010101000";
                when x"66" => data <= "0100000000";
                when x"67" => data <= "0100000000";
                when x"68" => data <= "0101011111";
                when x"69" => data <= "0010101000";
                when x"6A" => data <= "1111111000";
                when x"6B" => data <= "0100000000";
                when x"6C" => data <= "1001111111";
                when x"6D" => data <= "1000010101";
                when x"6E" => data <= "1111010111";
                when x"6F" => data <= "0111111011";
                when x"70" => data <= "1001111111";
                when x"71" => data <= "0111001110";
                when x"72" => data <= "1010101011";
                when x"73" => data <= "1110111101";
                when x"74" => data <= "0111111011";
                when x"75" => data <= "0101110000";
                when x"76" => data <= "1001111111";
                when x"77" => data <= "1111010111";
                when x"78" => data <= "0111111011";
                when x"79" => data <= "1001111111";
                when x"7A" => data <= "0000001100";
                when x"7B" => data <= "0101110000";
                when x"7C" => data <= "1000100000";
                when x"7D" => data <= "1001111111";
                when x"7E" => data <= "1001111111";
                when x"7F" => data <= "1110111101";
                when x"80" => data <= "1111010111";
                when x"81" => data <= "1110111101";
                when x"82" => data <= "0111111011";
                when x"83" => data <= "0011101101";
                when x"84" => data <= "0101000101";
                when x"85" => data <= "0111111011";
                when x"86" => data <= "0100101111";
                when x"87" => data <= "0100101111";
                when x"88" => data <= "0111111011";
                when x"89" => data <= "1110001000";
                when x"8A" => data <= "0100101111";
                when x"8B" => data <= "1111010111";
                when x"8C" => data <= "1001111111";
                when x"8D" => data <= "1111010111";
                when x"8E" => data <= "0111111011";
                when x"8F" => data <= "1001111111";
                when x"90" => data <= "0111111011";
                when x"91" => data <= "1110111101";
                when x"92" => data <= "1000100000";
                when x"93" => data <= "0001010011";
                when x"94" => data <= "1001111111";
                when x"95" => data <= "0111001110";
                when x"96" => data <= "0111111011";
                when x"97" => data <= "0111111011";
                when x"98" => data <= "1001111111";
                when x"99" => data <= "0111111011";
                when x"9A" => data <= "0111111011";
                when x"9B" => data <= "0111001110";
                when x"9C" => data <= "0000001100";
                when x"9D" => data <= "0101000101";
                when x"9E" => data <= "1110111101";
                when x"9F" => data <= "0111111011";
                when x"A0" => data <= "1000010101";
                when x"A1" => data <= "1110001000";
                when x"A2" => data <= "1101011100";
                when x"A3" => data <= "1001111111";
                when x"A4" => data <= "0011011000";
                when x"A5" => data <= "1110001000";
                when x"A6" => data <= "1110111101";
                when x"A7" => data <= "0101000101";
                when x"A8" => data <= "0100101111";
                when x"A9" => data <= "0111001110";
                when x"AA" => data <= "1110111101";
                when x"AB" => data <= "0110000110";
                when x"AC" => data <= "1100010100";
                when x"AD" => data <= "0101010010";
                when x"AE" => data <= "1111000000";
                when x"AF" => data <= "1000000010";
                when x"B0" => data <= "0110000110";
                when x"B1" => data <= "1111110101";
                when x"B2" => data <= "1111000000";
                when x"B3" => data <= "0001000100";
                when x"B4" => data <= "0100111000";
                when x"B5" => data <= "0001000100";
                when x"B6" => data <= "1000110111";
                when x"B7" => data <= "1111110101";
                when x"B8" => data <= "1011010110";
                when x"B9" => data <= "0100001101";
                when x"BA" => data <= "0001000100";
                when x"BB" => data <= "0001000100";
                when x"BC" => data <= "0100001101";
                when x"BD" => data <= "1111000000";
                when x"BE" => data <= "0100111000";
                when x"BF" => data <= "1000110111";
                when x"C0" => data <= "1011100011";
                when x"C1" => data <= "1111000000";
                when x"C2" => data <= "0101010010";
                when x"C3" => data <= "1111000000";
                when x"C4" => data <= "1111110101";
                when x"C5" => data <= "0001000100";
                when x"C6" => data <= "0101010010";
                when x"C7" => data <= "1001011101";
                when x"C8" => data <= "0001000100";
                when x"C9" => data <= "1000000010";
                when x"CA" => data <= "0001000100";
                when x"CB" => data <= "0011111010";
                when x"CC" => data <= "0100001101";
                when x"CD" => data <= "0001000100";
                when x"CE" => data <= "0101100111";
                when x"CF" => data <= "1100010100";
                when x"D0" => data <= "0101010010";
                when x"D1" => data <= "0110000110";
                when x"D2" => data <= "0010100101";
                when x"D3" => data <= "1111011010";
                when x"D4" => data <= "1111011010";
                when x"D5" => data <= "1111011010";
                when x"D6" => data <= "1001110010";
                when x"D7" => data <= "0101001000";
                when x"D8" => data <= "0000000001";
                when x"D9" => data <= "1111101111";
                when x"DA" => data <= "1111011010";
                when x"DB" => data <= "1111011010";
                when x"DC" => data <= "1111101111";
                when x"DD" => data <= "1111011010";
                when x"DE" => data <= "1011001100";
                when x"DF" => data <= "1000011000";
                when x"E0" => data <= "0010111111";
                when x"E1" => data <= "1111101111";
                when x"E2" => data <= "1011111001";
                when x"E3" => data <= "1111101111";
                when x"E4" => data <= "1111011010";
                when x"E5" => data <= "1111011010";
                when x"E6" => data <= "1111011010";
                when x"E7" => data <= "1001110010";
                when x"E8" => data <= "0000000001";
                when x"E9" => data <= "1100111011";
                when x"EA" => data <= "1111011010";
                when x"EB" => data <= "1111011010";
                when x"EC" => data <= "1111101111";
                when x"ED" => data <= "0000000001";
                when x"EE" => data <= "1111101111";
                when x"EF" => data <= "0010001010";
                when x"F0" => data <= "1111011010";
                when x"F1" => data <= "1000101101";
                when x"F2" => data <= "1111101111";
                when x"F3" => data <= "0110011100";
                when x"F4" => data <= "1111011010";
                when x"F5" => data <= "0010001010";
                when x"F6" => data <= "0000000001";
                when x"F7" => data <= "1111011010";
                when x"F8" => data <= "1011111001";
                when x"F9" => data <= "1111011010";
                when x"FA" => data <= "0000000001";
                when x"FB" => data <= "0110101001";
                when x"FC" => data <= "0101111101";
                when x"FD" => data <= "1111011010";
                when x"FE" => data <= "1111011010";
                when x"FF" => data <= "0100100010";
                when x"100" => data <= "0010111111";
                when x"101" => data <= "1001000111";
                when x"102" => data <= "1111011010";
                when x"103" => data <= "1111011010";
                when x"104" => data <= "1000011000";
                when x"105" => data <= "0110011100";
                when x"106" => data <= "1111011010";
                when x"107" => data <= "0100010111";
                when x"108" => data <= "1000101101";
                when x"109" => data <= "0000000001";
                when x"10A" => data <= "0000000001";
                when x"10B" => data <= "0110101001";
                when x"10C" => data <= "1100111011";
                when x"10D" => data <= "1100111011";
                when x"10E" => data <= "0010001010";
                when x"10F" => data <= "1111101111";
                when x"110" => data <= "1000101101";
                when x"111" => data <= "1100001110";
                when x"112" => data <= "1000101101";
                when x"113" => data <= "1111011010";
                when x"114" => data <= "1111011010";
                when x"115" => data <= "1111011010";
                when x"116" => data <= "0000000001";
                when x"117" => data <= "0111111101";
                when x"118" => data <= "0010000001";
                when x"119" => data <= "0000001010";
                when x"11A" => data <= "0111111101";
                when x"11B" => data <= "1101011010";
                when x"11C" => data <= "1101011010";
                when x"11D" => data <= "0110100010";
                when x"11E" => data <= "1010101101";
                when x"11F" => data <= "1110111011";
                when x"120" => data <= "0000111111";
                when x"121" => data <= "1101011010";
                when x"122" => data <= "0111001000";
                when x"123" => data <= "1010101101";
                when x"124" => data <= "0000111111";
                when x"125" => data <= "1010101101";
                when x"126" => data <= "1010101101";
                when x"127" => data <= "1110111011";
                when x"128" => data <= "1010011000";
                when x"129" => data <= "0111001000";
                when x"12A" => data <= "0100101001";
                when x"12B" => data <= "0111001000";
                when x"12C" => data <= "1110001110";
                when x"12D" => data <= "1100110000";
                when x"12E" => data <= "0100101001";
                when x"12F" => data <= "0111001000";
                when x"130" => data <= "0000001010";
                when x"131" => data <= "1010011000";
                when x"132" => data <= "0111111101";
                when x"133" => data <= "1101011010";
                when x"134" => data <= "0011101011";
                when x"135" => data <= "1010101101";
                when x"136" => data <= "0111111101";
                when x"137" => data <= "1110111011";
                when x"138" => data <= "1010101101";
                when x"139" => data <= "0100101001";
                when x"13A" => data <= "1110111011";
                when x"13B" => data <= "1110111011";
                when x"13C" => data <= "0001010101";
                when x"13D" => data <= "1111111110";
                when x"13E" => data <= "1011101000";
                when x"13F" => data <= "1111111110";
                when x"140" => data <= "0000010000";
                when x"141" => data <= "0000100101";
                when x"142" => data <= "1111111110";
                when x"143" => data <= "0001001111";
                when x"144" => data <= "0111100111";
                when x"145" => data <= "0111100111";
                when x"146" => data <= "0100000110";
                when x"147" => data <= "0100110011";
                when x"148" => data <= "0000100101";
                when x"149" => data <= "1000001001";
                when x"14A" => data <= "1000001001";
                when x"14B" => data <= "0000100101";
                when x"14C" => data <= "0100000110";
                when x"14D" => data <= "0000100101";
                when x"14E" => data <= "1010000010";
                when x"14F" => data <= "0111100111";
                when x"150" => data <= "0000010000";
                when x"151" => data <= "0111010010";
                when x"152" => data <= "0100000110";
                when x"153" => data <= "1111111110";
                when x"154" => data <= "1111111110";
                when x"155" => data <= "0000100101";
                when x"156" => data <= "0000100101";
                when x"157" => data <= "0111010010";
                when x"158" => data <= "1111111110";
                when x"159" => data <= "0110001101";
                when x"15A" => data <= "1011101000";
                when x"15B" => data <= "0000010000";
                when x"15C" => data <= "0000100101";
                when x"15D" => data <= "0000100101";
                when x"15E" => data <= "1111111110";
                when x"15F" => data <= "0001111010";
                when x"160" => data <= "1111111110";
                when x"161" => data <= "0100000110";
                when x"162" => data <= "1111111110";
                when x"163" => data <= "0000100101";
                when x"164" => data <= "0111100111";
                when x"165" => data <= "0111100111";
                when x"166" => data <= "1111111110";
                when x"167" => data <= "1111111110";
                when x"168" => data <= "0000100101";
                when x"169" => data <= "0000100101";
                when x"16A" => data <= "0100000110";
                when x"16B" => data <= "1000111100";
                when x"16C" => data <= "0011000100";
                when x"16D" => data <= "1000001001";
                when x"16E" => data <= "1111111110";
                when x"16F" => data <= "1111111110";
                when x"170" => data <= "0000010000";
                when x"171" => data <= "0000100101";
                when x"172" => data <= "0111010010";
                when x"173" => data <= "0000100101";
                when x"174" => data <= "1111111110";
                when x"175" => data <= "1000001001";
                when x"176" => data <= "0000100101";
                when x"177" => data <= "1111111110";
                when x"178" => data <= "1111111110";
                when x"179" => data <= "0000100101";
                when x"17A" => data <= "0011000100";
                when x"17B" => data <= "0000010000";
                when x"17C" => data <= "0100110011";
                when x"17D" => data <= "1111111110";
                when x"17E" => data <= "0000100101";
                when x"17F" => data <= "0000010000";
                when x"180" => data <= "0110011010";
                when x"181" => data <= "0100100100";
                when x"182" => data <= "1011111111";
                when x"183" => data <= "1011111111";
                when x"184" => data <= "1011111111";
                when x"185" => data <= "1011111111";
                when x"186" => data <= "1011111111";
                when x"187" => data <= "0110101111";
                when x"188" => data <= "0110101111";
                when x"189" => data <= "1011111111";
                when x"18A" => data <= "1011111111";
                when x"18B" => data <= "1011111111";
                when x"18C" => data <= "0001011000";
                when x"18D" => data <= "1011111111";
                when x"18E" => data <= "1011111111";
                when x"18F" => data <= "1011111111";
                when x"190" => data <= "1011111111";
                when x"191" => data <= "0001101101";
                when x"192" => data <= "1001000001";
                when x"193" => data <= "1011111111";
                when x"194" => data <= "1011111111";
                when x"195" => data <= "0001101101";
                when x"196" => data <= "1011111111";
                when x"197" => data <= "1011111111";
                when x"198" => data <= "1011111111";
                when x"199" => data <= "1011111111";
                when x"19A" => data <= "1011111111";
                when x"19B" => data <= "1011111111";
                when x"19C" => data <= "1011111111";
                when x"19D" => data <= "1011111111";
                when x"19E" => data <= "1011111111";
                when x"19F" => data <= "1011111111";
                when x"1A0" => data <= "0010001100";
                when x"1A1" => data <= "1011111111";
                when x"1A2" => data <= "1011111111";
                when x"1A3" => data <= "1011111111";
                when x"1A4" => data <= "1011111111";
                when x"1A5" => data <= "1011111111";
                when x"1A6" => data <= "1011111111";
                when x"1A7" => data <= "1011111111";
                when x"1A8" => data <= "1011111111";
                when x"1A9" => data <= "0110101111";
                when x"1AA" => data <= "1011111111";
                when x"1AB" => data <= "1011111111";
                when x"1AC" => data <= "1011111111";
                when x"1AD" => data <= "1011111111";
                when x"1AE" => data <= "1011111111";
                when x"1AF" => data <= "1011111111";
                when x"1B0" => data <= "1100001000";
                when x"1B1" => data <= "1101010111";
                when x"1B2" => data <= "1011111111";
                when x"1B3" => data <= "0001011000";
                when x"1B4" => data <= "1011111111";
                when x"1B5" => data <= "1010100000";
                when x"1B6" => data <= "1110110110";
                when x"1B7" => data <= "0110011010";
                when x"1B8" => data <= "0010001100";
                when x"1B9" => data <= "0101111011";
                when x"1BA" => data <= "1011111111";
                when x"1BB" => data <= "1011111111";
                when x"1BC" => data <= "1011111111";
                when x"1BD" => data <= "1011111111";
                when x"1BE" => data <= "1011111111";
                when x"1BF" => data <= "1011111111";
                when x"1C0" => data <= "1011111111";
                when x"1C1" => data <= "1011111111";
                when x"1C2" => data <= "1011111111";
                when x"1C3" => data <= "1011111111";
                when x"1C4" => data <= "0100100100";
                when x"1C5" => data <= "0001101101";
                when x"1C6" => data <= "1011111111";
                when x"1C7" => data <= "1011001010";
                when x"1C8" => data <= "1011111111";
                when x"1C9" => data <= "1011111111";
                when x"1CA" => data <= "1101010111";
                when x"1CB" => data <= "1011111111";
                when x"1CC" => data <= "0110101111";
                when x"1CD" => data <= "0000000111";
                when x"1CE" => data <= "1011111111";
                when x"1CF" => data <= "1011111111";
                when x"1D0" => data <= "1011111111";
                when x"1D1" => data <= "0110101111";
                when x"1D2" => data <= "1011111111";
                when x"1D3" => data <= "1011111111";
                when x"1D4" => data <= "1011111111";
                when x"1D5" => data <= "1011111111";
                when x"1D6" => data <= "1011111111";
                when x"1D7" => data <= "1011111111";
                when x"1D8" => data <= "1011111111";
                when x"1D9" => data <= "1011111111";
                when x"1DA" => data <= "1011111111";
                when x"1DB" => data <= "0101111011";
                when x"1DC" => data <= "1011111111";
                when x"1DD" => data <= "1011111111";
                when x"1DE" => data <= "0110011010";
                when x"1DF" => data <= "0110101111";
                when x"1E0" => data <= "1011111111";
                when x"1E1" => data <= "1011111111";
                when x"1E2" => data <= "1011111111";
                when x"1E3" => data <= "1011111111";
                when x"1E4" => data <= "0110101111";
                when x"1E5" => data <= "1011111111";
                when x"1E6" => data <= "1011111111";
                when x"1E7" => data <= "1100111101";
                when x"1E8" => data <= "1011111111";
                when x"1E9" => data <= "1011111111";
                when x"1EA" => data <= "1011111111";
                when x"1EB" => data <= "1011111111";
                when x"1EC" => data <= "1011111111";
                when x"1ED" => data <= "1011111111";
                when x"1EE" => data <= "1011111111";
                when x"1EF" => data <= "1010100000";
                when x"1F0" => data <= "1011111111";
                when x"1F1" => data <= "1011111111";
                when x"1F2" => data <= "1011111111";
                when x"1F3" => data <= "1011111111";
                when x"1F4" => data <= "1011111111";
                when x"1F5" => data <= "0110101111";
                when x"1F6" => data <= "1011111111";
                when x"1F7" => data <= "1011111111";
                when x"1F8" => data <= "1011111111";
                when x"1F9" => data <= "0110101111";
                when x"1FA" => data <= "1101010111";
                when x"1FB" => data <= "1011111111";
                when x"1FC" => data <= "1011111111";
                when x"1FD" => data <= "1101111000";
                when x"1FE" => data <= "0110000000";
                when x"1FF" => data <= "0100001011";
                when x"200" => data <= "0110000000";
                when x"201" => data <= "0110000000";
                when x"202" => data <= "1000000100";
                when x"203" => data <= "0111011111";
                when x"204" => data <= "1000110001";
                when x"205" => data <= "1111110011";
                when x"206" => data <= "0001000010";
                when x"207" => data <= "0110000000";
                when x"208" => data <= "0000101000";
                when x"209" => data <= "0000101000";
                when x"20A" => data <= "0110000000";
                when x"20B" => data <= "0110000000";
                when x"20C" => data <= "1100100111";
                when x"20D" => data <= "0111011111";
                when x"20E" => data <= "1000000100";
                when x"20F" => data <= "0111011111";
                when x"210" => data <= "1000000100";
                when x"211" => data <= "0000101000";
                when x"212" => data <= "0101010100";
                when x"213" => data <= "1000000100";
                when x"214" => data <= "1011010000";
                when x"215" => data <= "1000000100";
                when x"216" => data <= "0111011111";
                when x"217" => data <= "1000110001";
                when x"218" => data <= "1001011011";
                when x"219" => data <= "0001000010";
                when x"21A" => data <= "0010100011";
                when x"21B" => data <= "1011010000";
                when x"21C" => data <= "0111011111";
                when x"21D" => data <= "0000101000";
                when x"21E" => data <= "1000000100";
                when x"21F" => data <= "0110000000";
                when x"220" => data <= "1000000100";
                when x"221" => data <= "1000000100";
                when x"222" => data <= "0110000000";
                when x"223" => data <= "1111110011";
                when x"224" => data <= "0000101000";
                when x"225" => data <= "0001000010";
                when x"226" => data <= "1000000100";
                when x"227" => data <= "1000000100";
                when x"228" => data <= "0000101000";
                when x"229" => data <= "0111011111";
                when x"22A" => data <= "0101010100";
                when x"22B" => data <= "0111011111";
                when x"22C" => data <= "0100001011";
                when x"22D" => data <= "1011010000";
                when x"22E" => data <= "0110000000";
                when x"22F" => data <= "1001011011";
                when x"230" => data <= "0110000000";
                when x"231" => data <= "0110000000";
                when x"232" => data <= "1000000100";
                when x"233" => data <= "0111011111";
                when x"234" => data <= "0110000000";
                when x"235" => data <= "0111011111";
                when x"236" => data <= "0110000000";
                when x"237" => data <= "1000000100";
                when x"238" => data <= "0001000010";
                when x"239" => data <= "0111011111";
                when x"23A" => data <= "1000000100";
                when x"23B" => data <= "1000000100";
                when x"23C" => data <= "1000000100";
                when x"23D" => data <= "0111011111";
                when x"23E" => data <= "0000101000";
                when x"23F" => data <= "1000000100";
                when x"240" => data <= "0000101000";
                when x"241" => data <= "1000000100";
                when x"242" => data <= "1111110110";
                when x"243" => data <= "1010111111";
                when x"244" => data <= "0111011010";
                when x"245" => data <= "0111101111";
                when x"246" => data <= "1010001010";
                when x"247" => data <= "1010111111";
                when x"248" => data <= "0000101101";
                when x"249" => data <= "0111011010";
                when x"24A" => data <= "1010111111";
                when x"24B" => data <= "0000101101";
                when x"24C" => data <= "1010111111";
                when x"24D" => data <= "0111011010";
                when x"24E" => data <= "0100111011";
                when x"24F" => data <= "0111101111";
                when x"250" => data <= "0000011000";
                when x"251" => data <= "1000110100";
                when x"252" => data <= "0000011000";
                when x"253" => data <= "1010001010";
                when x"254" => data <= "0000101101";
                when x"255" => data <= "0000101101";
                when x"256" => data <= "0111101111";
                when x"257" => data <= "0000101101";
                when x"258" => data <= "1111110110";
                when x"259" => data <= "1000000001";
                when x"25A" => data <= "1010111111";
                when x"25B" => data <= "0000101101";
                when x"25C" => data <= "1010111111";
                when x"25D" => data <= "1101111101";
                when x"25E" => data <= "0000101101";
                when x"25F" => data <= "1010111111";
                when x"260" => data <= "0000101101";
                when x"261" => data <= "0111101111";
                when x"262" => data <= "0000011000";
                when x"263" => data <= "0111011010";
                when x"264" => data <= "1000000001";
                when x"265" => data <= "1101111101";
                when x"266" => data <= "1010111111";
                when x"267" => data <= "1010111111";
                when x"268" => data <= "0111101111";
                when x"269" => data <= "1110011100";
                when x"26A" => data <= "1101111101";
                when x"26B" => data <= "0000101101";
                when x"26C" => data <= "0111101111";
                when x"26D" => data <= "0111101111";
                when x"26E" => data <= "0111011010";
                when x"26F" => data <= "0111101111";
                when x"270" => data <= "0100111011";
                when x"271" => data <= "1101111101";
                when x"272" => data <= "1101111101";
                when x"273" => data <= "1010111111";
                when x"274" => data <= "1010111111";
                when x"275" => data <= "1101111101";
                when x"276" => data <= "0111101111";
                when x"277" => data <= "0111011010";
                when x"278" => data <= "0000011000";
                when x"279" => data <= "0001000111";
                when x"27A" => data <= "0111101111";
                when x"27B" => data <= "0000101101";
                when x"27C" => data <= "0111101111";
                when x"27D" => data <= "1010111111";
                when x"27E" => data <= "0111101111";
                when x"27F" => data <= "1000000001";
                when x"280" => data <= "0100111011";
                when x"281" => data <= "0111101111";
                when x"282" => data <= "1010111111";
                when x"283" => data <= "0111101111";
                when x"284" => data <= "1000110100";
                when x"285" => data <= "1000000001";
                when x"286" => data <= "1101111101";
                when x"287" => data <= "1010001010";
                when x"288" => data <= "1101010010";
                when x"289" => data <= "1001110001";
                when x"28A" => data <= "0000000010";
                when x"28B" => data <= "0000000010";
                when x"28C" => data <= "0000000010";
                when x"28D" => data <= "1110000110";
                when x"28E" => data <= "0000000010";
                when x"28F" => data <= "0000000010";
                when x"290" => data <= "1001000100";
                when x"291" => data <= "0000000010";
                when x"292" => data <= "0000000010";
                when x"293" => data <= "0111110101";
                when x"294" => data <= "1011111010";
                when x"295" => data <= "1011111010";
                when x"296" => data <= "1001110001";
                when x"297" => data <= "1101010010";
                when x"298" => data <= "0111000000";
                when x"299" => data <= "1101010010";
                when x"29A" => data <= "1011111010";
                when x"29B" => data <= "0100010100";
                when x"29C" => data <= "0110101010";
                when x"29D" => data <= "1010100101";
                when x"29E" => data <= "1010100101";
                when x"29F" => data <= "0000000010";
                when x"2A0" => data <= "0100010100";
                when x"2A1" => data <= "1011111010";
                when x"2A2" => data <= "0111110101";
                when x"2A3" => data <= "0111000000";
                when x"2A4" => data <= "0000000010";
                when x"2A5" => data <= "0111000000";
                when x"2A6" => data <= "0111000000";
                when x"2A7" => data <= "1100001101";
                when x"2A8" => data <= "0000000010";
                when x"2A9" => data <= "1010100101";
                when x"2AA" => data <= "0110011111";
                when x"2AB" => data <= "0000000010";
                when x"2AC" => data <= "0000000010";
                when x"2AD" => data <= "0011010110";
                when x"2AE" => data <= "0100010100";
                when x"2AF" => data <= "1110000110";
                when x"2B0" => data <= "0000000010";
                when x"2B1" => data <= "1001110001";
                when x"2B2" => data <= "0110101010";
                when x"2B3" => data <= "0110011111";
                when x"2B4" => data <= "1001000100";
                when x"2B5" => data <= "1111011001";
                when x"2B6" => data <= "1011111010";
                when x"2B7" => data <= "1111111011";
                when x"2B8" => data <= "1111111011";
                when x"2B9" => data <= "0110001000";
                when x"2BA" => data <= "1111111011";
                when x"2BB" => data <= "1111111011";
                when x"2BC" => data <= "1111111011";
                when x"2BD" => data <= "0111010111";
                when x"2BE" => data <= "1000111001";
                when x"2BF" => data <= "0000100000";
                when x"2C0" => data <= "1000111001";
                when x"2C1" => data <= "0000100000";
                when x"2C2" => data <= "1011011000";
                when x"2C3" => data <= "0110001000";
                when x"2C4" => data <= "0000100000";
                when x"2C5" => data <= "1000111001";
                when x"2C6" => data <= "1011011000";
                when x"2C7" => data <= "0000010101";
                when x"2C8" => data <= "1111111011";
                when x"2C9" => data <= "0000100000";
                when x"2CA" => data <= "0110001000";
                when x"2CB" => data <= "1111111011";
                when x"2CC" => data <= "0111010111";
                when x"2CD" => data <= "1111111011";
                when x"2CE" => data <= "1111111011";
                when x"2CF" => data <= "1011101101";
                when x"2D0" => data <= "0110001000";
                when x"2D1" => data <= "0100000011";
                when x"2D2" => data <= "1011011000";
                when x"2D3" => data <= "0100000011";
                when x"2D4" => data <= "1111111011";
                when x"2D5" => data <= "0000100000";
                when x"2D6" => data <= "0010101011";
                when x"2D7" => data <= "1111111011";
                when x"2D8" => data <= "0000100000";
                when x"2D9" => data <= "1111111011";
                when x"2DA" => data <= "0000100000";
                when x"2DB" => data <= "0001111111";
                when x"2DC" => data <= "0000100000";
                when x"2DD" => data <= "0000010101";
                when x"2DE" => data <= "1111111011";
                when x"2DF" => data <= "1111111011";
                when x"2E0" => data <= "1111111011";
                when x"2E1" => data <= "1111111011";
                when x"2E2" => data <= "1111111011";
                when x"2E3" => data <= "0000100000";
                when x"2E4" => data <= "0000100000";
                when x"2E5" => data <= "0000100000";
                when x"2E6" => data <= "0000100000";
                when x"2E7" => data <= "0110001000";
                when x"2E8" => data <= "0000100000";
                when x"2E9" => data <= "0110001000";
                when x"2EA" => data <= "0001001010";
                when x"2EB" => data <= "1111111011";
                when x"2EC" => data <= "0000100000";
                when x"2ED" => data <= "0111010111";
                when x"2EE" => data <= "1111111011";
                when x"2EF" => data <= "1111111011";
                when x"2F0" => data <= "1011101101";
                when x"2F1" => data <= "1111111011";
                when x"2F2" => data <= "0111100010";
                when x"2F3" => data <= "0000100000";
                when x"2F4" => data <= "1111111011";
                when x"2F5" => data <= "0000100000";
                when x"2F6" => data <= "1111111011";
                when x"2F7" => data <= "1111111011";
                when x"2F8" => data <= "1111111011";
                when x"2F9" => data <= "1111111011";
                when x"2FA" => data <= "0000100000";
                when x"2FB" => data <= "0010101011";
                when x"2FC" => data <= "1111111011";
                when x"2FD" => data <= "0000100000";
                when x"2FE" => data <= "1111111011";
                when x"2FF" => data <= "1111111011";
                when x"300" => data <= "0000100000";
                when x"301" => data <= "1100011010";
                when x"302" => data <= "1111111011";
                when x"303" => data <= "0000100000";
                when x"304" => data <= "1111111011";
                when x"305" => data <= "1111111011";
                when x"306" => data <= "1111111011";
                when x"307" => data <= "0000100000";
                when x"308" => data <= "0000100000";
                when x"309" => data <= "1011011000";
                when x"30A" => data <= "1111111011";
                when x"30B" => data <= "1100101111";
                when x"30C" => data <= "1111111011";
                when x"30D" => data <= "1000111001";
                when x"30E" => data <= "1111111011";
                when x"30F" => data <= "1111111011";
                when x"310" => data <= "1111111011";
                when x"311" => data <= "1011000010";
                when x"312" => data <= "0001010000";
                when x"313" => data <= "1000010110";
                when x"314" => data <= "1111010100";
                when x"315" => data <= "1011110111";
                when x"316" => data <= "1111010100";
                when x"317" => data <= "0101000110";
                when x"318" => data <= "1100000000";
                when x"319" => data <= "0101110011";
                when x"31A" => data <= "1011110111";
                when x"31B" => data <= "1001001001";
                when x"31C" => data <= "1011110111";
                when x"31D" => data <= "1110001011";
                when x"31E" => data <= "1010101000";
                when x"31F" => data <= "1000010110";
                when x"320" => data <= "1000100011";
                when x"321" => data <= "0001010000";
                when x"322" => data <= "0001010000";
                when x"323" => data <= "0001010000";
                when x"324" => data <= "1010101000";
                when x"325" => data <= "0001010000";
                when x"326" => data <= "0001010000";
                when x"327" => data <= "1100000000";
                when x"328" => data <= "0110100111";
                when x"329" => data <= "1101011111";
                when x"32A" => data <= "1101011111";
                when x"32B" => data <= "0010000100";
                when x"32C" => data <= "0110100111";
                when x"32D" => data <= "1100000000";
                when x"32E" => data <= "0001100101";
                when x"32F" => data <= "1010101000";
                when x"330" => data <= "1011110111";
                when x"331" => data <= "0001010000";
                when x"332" => data <= "0110100111";
                when x"333" => data <= "1011110111";
                when x"334" => data <= "0010000100";
                when x"335" => data <= "1110111110";
                when x"336" => data <= "0110100111";
                when x"337" => data <= "1010101000";
                when x"338" => data <= "1010101000";
                when x"339" => data <= "1100000000";
                when x"33A" => data <= "1011110111";
                when x"33B" => data <= "1101011111";
                when x"33C" => data <= "1011110111";
                when x"33D" => data <= "1100110101";
                when x"33E" => data <= "1101011111";
                when x"33F" => data <= "0101000110";
                when x"340" => data <= "0010000100";
                when x"341" => data <= "1000100011";
                when x"342" => data <= "1011110111";
                when x"343" => data <= "1001000010";
                when x"344" => data <= "0000000100";
                when x"345" => data <= "0000000100";
                when x"346" => data <= "1111011111";
                when x"347" => data <= "0000000100";
                when x"348" => data <= "1001000010";
                when x"349" => data <= "1111011111";
                when x"34A" => data <= "1111011111";
                when x"34B" => data <= "1001110111";
                when x"34C" => data <= "1111011111";
                when x"34D" => data <= "0111000110";
                when x"34E" => data <= "1111011111";
                when x"34F" => data <= "0000000100";
                when x"350" => data <= "0000000100";
                when x"351" => data <= "0111000110";
                when x"352" => data <= "1001110111";
                when x"353" => data <= "0000000100";
                when x"354" => data <= "0000000100";
                when x"355" => data <= "0000000100";
                when x"356" => data <= "1000101000";
                when x"357" => data <= "0000000100";
                when x"358" => data <= "0000000100";
                when x"359" => data <= "1111011111";
                when x"35A" => data <= "0000000100";
                when x"35B" => data <= "1001000010";
                when x"35C" => data <= "1111011111";
                when x"35D" => data <= "0000000100";
                when x"35E" => data <= "0000000100";
                when x"35F" => data <= "0000000100";
                when x"360" => data <= "1000101000";
                when x"361" => data <= "0000000100";
                when x"362" => data <= "0000000100";
                when x"363" => data <= "1110110101";
                when x"364" => data <= "1001000010";
                when x"365" => data <= "1110000000";
                when x"366" => data <= "0000000100";
                when x"367" => data <= "0000000100";
                when x"368" => data <= "0000000100";
                when x"369" => data <= "1111011111";
                when x"36A" => data <= "1111011111";
                when x"36B" => data <= "1111011111";
                when x"36C" => data <= "0000000100";
                when x"36D" => data <= "0111000110";
                when x"36E" => data <= "0100010010";
                when x"36F" => data <= "1001000010";
                when x"370" => data <= "0000000100";
                when x"371" => data <= "1111101010";
                when x"372" => data <= "0010111010";
                when x"373" => data <= "1001110111";
                when x"374" => data <= "1110000000";
                when x"375" => data <= "1101010100";
                when x"376" => data <= "0000000100";
                when x"377" => data <= "0000000100";
                when x"378" => data <= "0100010010";
                when x"379" => data <= "1111011111";
                when x"37A" => data <= "0000000100";
                when x"37B" => data <= "1111011111";
                when x"37C" => data <= "0000000100";
                when x"37D" => data <= "0000000100";
                when x"37E" => data <= "1111011111";
                when x"37F" => data <= "0000000100";
                when x"380" => data <= "1000101000";
                when x"381" => data <= "0000000100";
                when x"382" => data <= "0011100101";
                when x"383" => data <= "0000000100";
                when x"384" => data <= "1001000010";
                when x"385" => data <= "0000000100";
                when x"386" => data <= "1111011111";
                when x"387" => data <= "0000000100";
                when x"388" => data <= "0100100111";
                when x"389" => data <= "0000000100";
                when x"38A" => data <= "0000000100";
                when x"38B" => data <= "1001110111";
                when x"38C" => data <= "0100010010";
                when x"38D" => data <= "0000000100";
                when x"38E" => data <= "1001110111";
                when x"38F" => data <= "1110000000";
                when x"390" => data <= "1001110111";
                when x"391" => data <= "1111011111";
                when x"392" => data <= "0000000100";
                when x"393" => data <= "1110000000";
                when x"394" => data <= "0000000100";
                when x"395" => data <= "1001110111";
                when x"396" => data <= "0000000100";
                when x"397" => data <= "1000101000";
                when x"398" => data <= "1111011111";
                when x"399" => data <= "1000011101";
                when x"39A" => data <= "1001000010";
                when x"39B" => data <= "0000000100";
                when x"39C" => data <= "0000000100";
                when x"39D" => data <= "0000000100";
                when x"39E" => data <= "0110101100";
                when x"39F" => data <= "0011111111";
                when x"3A0" => data <= "1001011000";
                when x"3A1" => data <= "0011111111";
                when x"3A2" => data <= "0100001000";
                when x"3A3" => data <= "0100001000";
                when x"3A4" => data <= "0011001010";
                when x"3A5" => data <= "0100111101";
                when x"3A6" => data <= "0000101011";
                when x"3A7" => data <= "1001011000";
                when x"3A8" => data <= "0011111111";
                when x"3A9" => data <= "1110101111";
                when x"3AA" => data <= "0100001000";
                when x"3AB" => data <= "1110011010";
                when x"3AC" => data <= "0100001000";
                when x"3AD" => data <= "0100001000";
                when x"3AE" => data <= "1001011000";
                when x"3AF" => data <= "1110011010";
                when x"3B0" => data <= "1001011000";
                when x"3B1" => data <= "0101100010";
                when x"3B2" => data <= "1110101111";
                when x"3B3" => data <= "0100001000";
                when x"3B4" => data <= "1010111001";
                when x"3B5" => data <= "1001011000";
                when x"3B6" => data <= "0010100000";
                when x"3B7" => data <= "1110101111";
                when x"3B8" => data <= "1110101111";
                when x"3B9" => data <= "1101111011";
                when x"3BA" => data <= "1101111011";
                when x"3BB" => data <= "0100111101";
                when x"3BC" => data <= "0101010111";
                when x"3BD" => data <= "0011111111";
                when x"3BE" => data <= "1001011000";
                when x"3BF" => data <= "1110101111";
                when x"3C0" => data <= "0011111111";
                when x"3C1" => data <= "1111110000";
                when x"3C2" => data <= "0011111111";
                when x"3C3" => data <= "0100111101";
                when x"3C4" => data <= "1101111011";
                when x"3C5" => data <= "0100001000";
                when x"3C6" => data <= "1101111011";
                when x"3C7" => data <= "0100001000";
                when x"3C8" => data <= "0011001010";
                when x"3C9" => data <= "1110101111";
                when x"3CA" => data <= "0011111111";
                when x"3CB" => data <= "0101010111";
                when x"3CC" => data <= "0100001000";
                when x"3CD" => data <= "0011001010";
                when x"3CE" => data <= "0100001000";
                when x"3CF" => data <= "1101111011";
                when x"3D0" => data <= "1011010011";
                when x"3D1" => data <= "0011111111";
                when x"3D2" => data <= "0100001000";
                when x"3D3" => data <= "0001000001";
                when x"3D4" => data <= "0011001010";
                when x"3D5" => data <= "0011001010";
                when x"3D6" => data <= "1000000111";
                when x"3D7" => data <= "0100111101";
                when x"3D8" => data <= "1110101111";
                when x"3D9" => data <= "0101000000";
                when x"3DA" => data <= "1000010000";
                when x"3DB" => data <= "0111111110";
                when x"3DC" => data <= "1000010000";
                when x"3DD" => data <= "1111010010";
                when x"3DE" => data <= "0101000000";
                when x"3DF" => data <= "1110111000";
                when x"3E0" => data <= "1111010010";
                when x"3E1" => data <= "1000010000";
                when x"3E2" => data <= "1100000110";
                when x"3E3" => data <= "0101000000";
                when x"3E4" => data <= "1110111000";
                when x"3E5" => data <= "1000010000";
                when x"3E6" => data <= "0101110101";
                when x"3E7" => data <= "1110111000";
                when x"3E8" => data <= "0111111110";
                when x"3E9" => data <= "1000100101";
                when x"3EA" => data <= "1011110001";
                when x"3EB" => data <= "0010000010";
                when x"3EC" => data <= "1101011001";
                when x"3ED" => data <= "0101000000";
                when x"3EE" => data <= "1000010000";
                when x"3EF" => data <= "0101110101";
                when x"3F0" => data <= "0101000000";
                when x"3F1" => data <= "0000001001";
                when x"3F2" => data <= "1000010000";
                when x"3F3" => data <= "1000010000";
                when x"3F4" => data <= "0101110101";
                when x"3F5" => data <= "0101000000";
                when x"3F6" => data <= "1111010010";
                when x"3F7" => data <= "1001111010";
                when x"3F8" => data <= "1110111000";
                when x"3F9" => data <= "1000010000";
                when x"3FA" => data <= "1111100111";
                when x"3FB" => data <= "1111010010";
                when x"3FC" => data <= "1000100101";
                when x"3FD" => data <= "0101000000";
                when x"3FE" => data <= "1000010000";
                when x"3FF" => data <= "1010101110";
                when x"400" => data <= "1111010010";
                when x"401" => data <= "1111010010";
                when x"402" => data <= "0001010110";
                when x"403" => data <= "0101000000";
                when x"404" => data <= "0010000010";
                when x"405" => data <= "0111001011";
                when x"406" => data <= "1000010000";
                when x"407" => data <= "0101110101";
                when x"408" => data <= "0101110101";
                when x"409" => data <= "0101110101";
                when x"40A" => data <= "1110111000";
                when x"40B" => data <= "0111001011";
                when x"40C" => data <= "1000010000";
                when x"40D" => data <= "0101000000";
                when x"40E" => data <= "0010000010";
                when x"40F" => data <= "0101110101";
                when x"410" => data <= "0101110101";
                when x"411" => data <= "0010000010";
                when x"412" => data <= "1010101110";
                when x"413" => data <= "1000100101";
                when x"414" => data <= "0101110101";
                when x"415" => data <= "0101110101";
                when x"416" => data <= "0101000000";
                when x"417" => data <= "0001010110";
                when x"418" => data <= "1000010000";
                when x"419" => data <= "1000100101";
                when x"41A" => data <= "1111111101";
                when x"41B" => data <= "0011110010";
                when x"41C" => data <= "0000010011";
                when x"41D" => data <= "1111001000";
                when x"41E" => data <= "0101011010";
                when x"41F" => data <= "1000111111";
                when x"420" => data <= "1011011110";
                when x"421" => data <= "1111111101";
                when x"422" => data <= "1111111101";
                when x"423" => data <= "0100000101";
                when x"424" => data <= "1110010111";
                when x"425" => data <= "1000111111";
                when x"426" => data <= "0101101111";
                when x"427" => data <= "1000001010";
                when x"428" => data <= "1011011110";
                when x"429" => data <= "0100000101";
                when x"42A" => data <= "1000001010";
                when x"42B" => data <= "1001010101";
                when x"42C" => data <= "1111001000";
                when x"42D" => data <= "1111111101";
                when x"42E" => data <= "1111001000";
                when x"42F" => data <= "1111111101";
                when x"430" => data <= "1011101011";
                when x"431" => data <= "0010011000";
                when x"432" => data <= "1111111101";
                when x"433" => data <= "1111111101";
                when x"434" => data <= "1011011110";
                when x"435" => data <= "0111010001";
                when x"436" => data <= "0100000101";
                when x"437" => data <= "1111111101";
                when x"438" => data <= "0001001100";
                when x"439" => data <= "1111111101";
                when x"43A" => data <= "0100000101";
                when x"43B" => data <= "1111111101";
                when x"43C" => data <= "1110010111";
                when x"43D" => data <= "1111111101";
                when x"43E" => data <= "1111111101";
                when x"43F" => data <= "1000111111";
                when x"440" => data <= "1111111101";
                when x"441" => data <= "1001010101";
                when x"442" => data <= "0101101111";
                when x"443" => data <= "1000001010";
                when x"444" => data <= "1000111111";
                when x"445" => data <= "1111111101";
                when x"446" => data <= "0100000101";
                when x"447" => data <= "0010101101";
                when x"448" => data <= "0100000101";
                when x"449" => data <= "1001100000";
                when x"44A" => data <= "1111111101";
                when x"44B" => data <= "1111111101";
                when x"44C" => data <= "1100111111";
                when x"44D" => data <= "1010100010";
                when x"44E" => data <= "1010010111";
                when x"44F" => data <= "1111011110";
                when x"450" => data <= "1100111111";
                when x"451" => data <= "1011111101";
                when x"452" => data <= "0010111011";
                when x"453" => data <= "1111011110";
                when x"454" => data <= "0110101101";
                when x"455" => data <= "0111000111";
                when x"456" => data <= "1100111111";
                when x"457" => data <= "0000000101";
                when x"458" => data <= "1011111101";
                when x"459" => data <= "0110101101";
                when x"45A" => data <= "1100111111";
                when x"45B" => data <= "0000000101";
                when x"45C" => data <= "1000011100";
                when x"45D" => data <= "1011111101";
                when x"45E" => data <= "1011111101";
                when x"45F" => data <= "0110101101";
                when x"460" => data <= "1110110100";
                when x"461" => data <= "0110101101";
                when x"462" => data <= "0000000101";
                when x"463" => data <= "0000000101";
                when x"464" => data <= "1011111101";
                when x"465" => data <= "1000101001";
                when x"466" => data <= "1111011110";
                when x"467" => data <= "1011111101";
                when x"468" => data <= "1100111111";
                when x"469" => data <= "0000000101";
                when x"46A" => data <= "1100111111";
                when x"46B" => data <= "0000000101";
                when x"46C" => data <= "0000000101";
                when x"46D" => data <= "0110101101";
                when x"46E" => data <= "1011001000";
                when x"46F" => data <= "0110011000";
                when x"470" => data <= "1100111111";
                when x"471" => data <= "1100111111";
                when x"472" => data <= "1011001000";
                when x"473" => data <= "0110101101";
                when x"474" => data <= "1010100010";
                when x"475" => data <= "0000000101";
                when x"476" => data <= "1000101001";
                when x"477" => data <= "1100111111";
                when x"478" => data <= "1111011110";
                when x"479" => data <= "0000000101";
                when x"47A" => data <= "1111011110";
                when x"47B" => data <= "0111000111";
                when x"47C" => data <= "1101010101";
                when x"47D" => data <= "0000000101";
                when x"47E" => data <= "0000000101";
                when x"47F" => data <= "1100111111";
                when x"480" => data <= "1100111111";
                when x"481" => data <= "1111101011";
                when x"482" => data <= "0000000101";
                when x"483" => data <= "1011111101";
                when x"484" => data <= "0000000101";
                when x"485" => data <= "0001011010";
                when x"486" => data <= "1011111101";
                when x"487" => data <= "0000000101";
                when x"488" => data <= "1011001000";
                when x"489" => data <= "0001000000";
                when x"48A" => data <= "0100001001";
                when x"48B" => data <= "0001000000";
                when x"48C" => data <= "1011010010";
                when x"48D" => data <= "0111011101";
                when x"48E" => data <= "1011100111";
                when x"48F" => data <= "0101010110";
                when x"490" => data <= "1101111010";
                when x"491" => data <= "0110000010";
                when x"492" => data <= "0001000000";
                when x"493" => data <= "0001000000";
                when x"494" => data <= "1011010010";
                when x"495" => data <= "0001000000";
                when x"496" => data <= "0001110101";
                when x"497" => data <= "0001000000";
                when x"498" => data <= "1011010010";
                when x"499" => data <= "0001000000";
                when x"49A" => data <= "0011001011";
                when x"49B" => data <= "1110101110";
                when x"49C" => data <= "1100010000";
                when x"49D" => data <= "0110000010";
                when x"49E" => data <= "1010111000";
                when x"49F" => data <= "0110000010";
                when x"4A0" => data <= "0001000000";
                when x"4A1" => data <= "0001000000";
                when x"4A2" => data <= "0010100001";
                when x"4A3" => data <= "1000110011";
                when x"4A4" => data <= "0001000000";
                when x"4A5" => data <= "1000110011";
                when x"4A6" => data <= "0001000000";
                when x"4A7" => data <= "0001000000";
                when x"4A8" => data <= "0001000000";
                when x"4A9" => data <= "0111101000";
                when x"4AA" => data <= "0001000000";
                when x"4AB" => data <= "1100010000";
                when x"4AC" => data <= "0001000000";
                when x"4AD" => data <= "0001000000";
                when x"4AE" => data <= "0100001001";
                when x"4AF" => data <= "0110000010";
                when x"4B0" => data <= "1111000100";
                when x"4B1" => data <= "0001000000";
                when x"4B2" => data <= "1011100111";
                when x"4B3" => data <= "0001000000";
                when x"4B4" => data <= "1011100111";
                when x"4B5" => data <= "0001000000";
                when x"4B6" => data <= "0001000000";
                when x"4B7" => data <= "0001000000";
                when x"4B8" => data <= "0001000000";
                when x"4B9" => data <= "0001000000";
                when x"4BA" => data <= "0001000000";
                when x"4BB" => data <= "0001000000";
                when x"4BC" => data <= "1010111000";
                when x"4BD" => data <= "0001000000";
                when x"4BE" => data <= "1011100111";
                when x"4BF" => data <= "1100100101";
                when x"4C0" => data <= "0001000000";
                when x"4C1" => data <= "0001000000";
                when x"4C2" => data <= "0001000000";
                when x"4C3" => data <= "1011100111";
                when x"4C4" => data <= "0000101010";
                when x"4C5" => data <= "0111101000";
                when x"4C6" => data <= "0001000000";
                when x"4C7" => data <= "0110110111";
                when x"4C8" => data <= "1011100111";
                when x"4C9" => data <= "0001000000";
                when x"4CA" => data <= "0001000000";
                when x"4CB" => data <= "0111101000";
                when x"4CC" => data <= "1001011001";
                when x"4CD" => data <= "1111000100";
                when x"4CE" => data <= "0111111111";
                when x"4CF" => data <= "0000001000";
                when x"4D0" => data <= "0111111111";
                when x"4D1" => data <= "0000001000";
                when x"4D2" => data <= "1000100100";
                when x"4D3" => data <= "1010101111";
                when x"4D4" => data <= "0111111111";
                when x"4D5" => data <= "1011000101";
                when x"4D6" => data <= "0000001000";
                when x"4D7" => data <= "0111111111";
                when x"4D8" => data <= "0111111111";
                when x"4D9" => data <= "0000001000";
                when x"4DA" => data <= "0111111111";
                when x"4DB" => data <= "0000001000";
                when x"4DC" => data <= "0000001000";
                when x"4DD" => data <= "0000001000";
                when x"4DE" => data <= "1001111011";
                when x"4DF" => data <= "0111111111";
                when x"4E0" => data <= "0111111111";
                when x"4E1" => data <= "1010101111";
                when x"4E2" => data <= "0111111111";
                when x"4E3" => data <= "0111001010";
                when x"4E4" => data <= "0111111111";
                when x"4E5" => data <= "0111111111";
                when x"4E6" => data <= "0000111101";
                when x"4E7" => data <= "0111111111";
                when x"4E8" => data <= "0000001000";
                when x"4E9" => data <= "0111111111";
                when x"4EA" => data <= "0111111111";
                when x"4EB" => data <= "0111111111";
                when x"4EC" => data <= "0111111111";
                when x"4ED" => data <= "0000001000";
                when x"4EE" => data <= "0111111111";
                when x"4EF" => data <= "0111111111";
                when x"4F0" => data <= "0111111111";
                when x"4F1" => data <= "0111111111";
                when x"4F2" => data <= "0111111111";
                when x"4F3" => data <= "0111111111";
                when x"4F4" => data <= "0111111111";
                when x"4F5" => data <= "1110111001";
                when x"4F6" => data <= "1010101111";
                when x"4F7" => data <= "0111111111";
                when x"4F8" => data <= "0111111111";
                when x"4F9" => data <= "0111111111";
                when x"4FA" => data <= "0000001000";
                when x"4FB" => data <= "0111111111";
                when x"4FC" => data <= "1000010001";
                when x"4FD" => data <= "0111111111";
                when x"4FE" => data <= "0000001000";
                when x"4FF" => data <= "0111111111";
                when x"500" => data <= "1001111011";
                when x"501" => data <= "0000001000";
                when x"502" => data <= "0000001000";
                when x"503" => data <= "1001111011";
                when x"504" => data <= "0000001000";
                when x"505" => data <= "0111111111";
                when x"506" => data <= "0111111111";
                when x"507" => data <= "1010101111";
                when x"508" => data <= "0000001000";
                when x"509" => data <= "0111111111";
                when x"50A" => data <= "0111111111";
                when x"50B" => data <= "0111111111";
                when x"50C" => data <= "1010101111";
                when x"50D" => data <= "0000001000";
                when x"50E" => data <= "0111111111";
                when x"50F" => data <= "0111111111";
                when x"510" => data <= "0111111111";
                when x"511" => data <= "0111111111";
                when x"512" => data <= "0111111111";
                when x"513" => data <= "0111111111";
                when x"514" => data <= "0111111111";
                when x"515" => data <= "1001111011";
                when x"516" => data <= "0000001000";
                when x"517" => data <= "1010101111";
                when x"518" => data <= "0111111111";
                when x"519" => data <= "0111111111";
                when x"51A" => data <= "0111111111";
                when x"51B" => data <= "0111111111";
                when x"51C" => data <= "0111111111";
                when x"51D" => data <= "0111111111";
                when x"51E" => data <= "0001010111";
                when x"51F" => data <= "0110100000";
                when x"520" => data <= "0111111111";
                when x"521" => data <= "0111111111";
                when x"522" => data <= "0111111111";
                when x"523" => data <= "0000001000";
                when x"524" => data <= "0111111111";
                when x"525" => data <= "0111111111";
                when x"526" => data <= "0111111111";
                when x"527" => data <= "1010101111";
                when x"528" => data <= "0111111111";
                when x"529" => data <= "0000001000";
                when x"52A" => data <= "0111111111";
                when x"52B" => data <= "0111111111";
                when x"52C" => data <= "0111111111";
                when x"52D" => data <= "0011101001";
                when x"52E" => data <= "0111111111";
                when x"52F" => data <= "0001010111";
                when x"530" => data <= "1001111011";
                when x"531" => data <= "0111001010";
                when x"532" => data <= "0000001000";
                when x"533" => data <= "0111111111";
                when x"534" => data <= "0111111111";
                when x"535" => data <= "0111111111";
                when x"536" => data <= "0000001000";
                when x"537" => data <= "0111111111";
                when x"538" => data <= "0111111111";
                when x"539" => data <= "0111111111";
                when x"53A" => data <= "0111111111";
                when x"53B" => data <= "0111111111";
                when x"53C" => data <= "0111111111";
                when x"53D" => data <= "0111111111";
                when x"53E" => data <= "0111111111";
                when x"53F" => data <= "0111111111";
                when x"540" => data <= "0000001000";
                when x"541" => data <= "0111111111";
                when x"542" => data <= "0111111111";
                when x"543" => data <= "0111111111";
                when x"544" => data <= "0111111111";
                when x"545" => data <= "0111111111";
                when x"546" => data <= "1010011010";
                when x"547" => data <= "0111111111";
                when x"548" => data <= "0111111111";
                when x"549" => data <= "0111111111";
                when x"54A" => data <= "0111111111";
                when x"54B" => data <= "0111111111";
                when x"54C" => data <= "0111111111";
                when x"54D" => data <= "0111111111";
                when x"54E" => data <= "0111111111";
                when x"54F" => data <= "0110100000";
                when x"550" => data <= "1000100100";
                when x"551" => data <= "1110111001";
                when x"552" => data <= "0111111111";
                when x"553" => data <= "0000001000";
                when x"554" => data <= "1010101111";
                when x"555" => data <= "0000001000";
                when x"556" => data <= "0111111111";
                when x"557" => data <= "0111111111";
                when x"558" => data <= "0111111111";
                when x"559" => data <= "0111111111";
                when x"55A" => data <= "0111111111";
                when x"55B" => data <= "0111111111";
                when x"55C" => data <= "0111111111";
                when x"55D" => data <= "0111111111";
                when x"55E" => data <= "0111111111";
                when x"55F" => data <= "0111111111";
                when x"560" => data <= "0111111111";
                when x"561" => data <= "0000001000";
                when x"562" => data <= "0000001000";
                when x"563" => data <= "0000001000";
                when x"564" => data <= "0111111111";
                when x"565" => data <= "0111111111";
                when x"566" => data <= "0111111111";
                when x"567" => data <= "0000001000";
                when x"568" => data <= "0000001000";
                when x"569" => data <= "0000001000";
                when x"56A" => data <= "0111111111";
                when x"56B" => data <= "0111111111";
                when x"56C" => data <= "0000001000";
                when x"56D" => data <= "0111111111";
                when x"56E" => data <= "0111111111";
                when x"56F" => data <= "0000001000";
                when x"570" => data <= "0111111111";
                when x"571" => data <= "0111111111";
                when x"572" => data <= "0000001000";
                when x"573" => data <= "0111111111";
                when x"574" => data <= "0000001000";
                when x"575" => data <= "0111111111";
                when x"576" => data <= "0111111111";
                when x"577" => data <= "0111111111";
                when x"578" => data <= "1001111011";
                when x"579" => data <= "0001010111";
                when x"57A" => data <= "0111111111";
                when x"57B" => data <= "0111111111";
                when x"57C" => data <= "0111111111";
                when x"57D" => data <= "0111111111";
                when x"57E" => data <= "0111111111";
                when x"57F" => data <= "1010011010";
                when x"580" => data <= "0111111111";
                when x"581" => data <= "0111111111";
                when x"582" => data <= "0000001000";
                when x"583" => data <= "0111111111";
                when x"584" => data <= "0000001000";
                when x"585" => data <= "0000001000";
                when x"586" => data <= "0111111111";
                when x"587" => data <= "0111111111";
                when x"588" => data <= "0111111111";
                when x"589" => data <= "0111111111";
                when x"58A" => data <= "0111111111";
                when x"58B" => data <= "0000010010";
                when x"58C" => data <= "0000010010";
                when x"58D" => data <= "1010000000";
                when x"58E" => data <= "1010000000";
                when x"58F" => data <= "0000100111";
                when x"590" => data <= "0000100111";
                when x"591" => data <= "1101110111";
                when x"592" => data <= "0110111010";
                when x"593" => data <= "1101110111";
                when x"594" => data <= "1101110111";
                when x"595" => data <= "1101110111";
                when x"596" => data <= "0111100101";
                when x"597" => data <= "0100000100";
                when x"598" => data <= "1010000000";
                when x"599" => data <= "1101110111";
                when x"59A" => data <= "1100101000";
                when x"59B" => data <= "1101110111";
                when x"59C" => data <= "1010000000";
                when x"59D" => data <= "0111100101";
                when x"59E" => data <= "0100000100";
                when x"59F" => data <= "0011110011";
                when x"5A0" => data <= "1111111100";
                when x"5A1" => data <= "0111100101";
                when x"5A2" => data <= "0100000100";
                when x"5A3" => data <= "0110111010";
                when x"5A4" => data <= "1011011111";
                when x"5A5" => data <= "0100000100";
                when x"5A6" => data <= "1101110111";
                when x"5A7" => data <= "1101110111";
                when x"5A8" => data <= "0100000100";
                when x"5A9" => data <= "1100011101";
                when x"5AA" => data <= "0011000110";
                when x"5AB" => data <= "1101110111";
                when x"5AC" => data <= "0010101100";
                when x"5AD" => data <= "1011011111";
                when x"5AE" => data <= "0100000100";
                when x"5AF" => data <= "1011011111";
                when x"5B0" => data <= "0100000100";
                when x"5B1" => data <= "1101110111";
                when x"5B2" => data <= "1100101000";
                when x"5B3" => data <= "0100000100";
                when x"5B4" => data <= "0111010000";
                when x"5B5" => data <= "1010000000";
                when x"5B6" => data <= "0111100101";
                when x"5B7" => data <= "1010000000";
                when x"5B8" => data <= "0100000100";
                when x"5B9" => data <= "0101011011";
                when x"5BA" => data <= "1010000000";
                when x"5BB" => data <= "0100000100";
                when x"5BC" => data <= "1100011101";
                when x"5BD" => data <= "1010000000";
                when x"5BE" => data <= "1101110111";
                when x"5BF" => data <= "1010000000";
                when x"5C0" => data <= "0100000100";
                when x"5C1" => data <= "1001010100";
                when x"5C2" => data <= "1010000000";
                when x"5C3" => data <= "1010000000";
                when x"5C4" => data <= "0010101100";
                when x"5C5" => data <= "0100000100";
                when x"5C6" => data <= "1101110111";
                when x"5C7" => data <= "1100011101";
                when x"5C8" => data <= "1101110111";
                when x"5C9" => data <= "1011011111";
                when x"5CA" => data <= "1101000010";
                when x"5CB" => data <= "0110111010";
                when x"5CC" => data <= "1101110111";
                when x"5CD" => data <= "0100000100";
                when x"5CE" => data <= "1000110101";
                when x"5CF" => data <= "1111110111";
                when x"5D0" => data <= "1000000000";
                when x"5D1" => data <= "1111110111";
                when x"5D2" => data <= "1111110111";
                when x"5D3" => data <= "1111110111";
                when x"5D4" => data <= "1000000000";
                when x"5D5" => data <= "1000000000";
                when x"5D6" => data <= "1000000000";
                when x"5D7" => data <= "1111110111";
                when x"5D8" => data <= "1000000000";
                when x"5D9" => data <= "1000000000";
                when x"5DA" => data <= "1000000000";
                when x"5DB" => data <= "1000000000";
                when x"5DC" => data <= "1000000000";
                when x"5DD" => data <= "1111110111";
                when x"5DE" => data <= "1000000000";
                when x"5DF" => data <= "1111110111";
                when x"5E0" => data <= "1010111110";
                when x"5E1" => data <= "1000000000";
                when x"5E2" => data <= "1000000000";
                when x"5E3" => data <= "0110000100";
                when x"5E4" => data <= "1000000000";
                when x"5E5" => data <= "1000000000";
                when x"5E6" => data <= "1000000000";
                when x"5E7" => data <= "1111110111";
                when x"5E8" => data <= "1000000000";
                when x"5E9" => data <= "1000110101";
                when x"5EA" => data <= "1000000000";
                when x"5EB" => data <= "1000000000";
                when x"5EC" => data <= "1000000000";
                when x"5ED" => data <= "1111110111";
                when x"5EE" => data <= "1111110111";
                when x"5EF" => data <= "1000000000";
                when x"5F0" => data <= "1111110111";
                when x"5F1" => data <= "1000000000";
                when x"5F2" => data <= "1000000000";
                when x"5F3" => data <= "1000000000";
                when x"5F4" => data <= "1111110111";
                when x"5F5" => data <= "1000000000";
                when x"5F6" => data <= "1000000000";
                when x"5F7" => data <= "1000000000";
                when x"5F8" => data <= "1000000000";
                when x"5F9" => data <= "1000110101";
                when x"5FA" => data <= "1000000000";
                when x"5FB" => data <= "1000000000";
                when x"5FC" => data <= "0111011011";
                when x"5FD" => data <= "1000000000";
                when x"5FE" => data <= "1000000000";
                when x"5FF" => data <= "0101100101";
                when x"600" => data <= "1111110111";
                when x"601" => data <= "1000000000";
                when x"602" => data <= "1000000000";
                when x"603" => data <= "1000000000";
                when x"604" => data <= "1111110111";
                when x"605" => data <= "1110101000";
                when x"606" => data <= "1000000000";
                when x"607" => data <= "1000000000";
                when x"608" => data <= "1111110111";
                when x"609" => data <= "1000000000";
                when x"60A" => data <= "1000000000";
                when x"60B" => data <= "1111110111";
                when x"60C" => data <= "1111110111";
                when x"60D" => data <= "1000000000";
                when x"60E" => data <= "1000000000";
                when x"60F" => data <= "1001011111";
                when x"610" => data <= "1111110111";
                when x"611" => data <= "1011100001";
                when x"612" => data <= "1000000000";
                when x"613" => data <= "1000000000";
                when x"614" => data <= "1111000010";
                when x"615" => data <= "0000101100";
                when x"616" => data <= "1000000000";
                when x"617" => data <= "1111110111";
                when x"618" => data <= "0101010000";
                when x"619" => data <= "1111110111";
                when x"61A" => data <= "1000000000";
                when x"61B" => data <= "1000000000";
                when x"61C" => data <= "1111110111";
                when x"61D" => data <= "1110101000";
                when x"61E" => data <= "1000000000";
                when x"61F" => data <= "1000000000";
                when x"620" => data <= "1000000000";
                when x"621" => data <= "1000000000";
                when x"622" => data <= "1000000000";
                when x"623" => data <= "1000000000";
                when x"624" => data <= "1000110101";
                when x"625" => data <= "1000000000";
                when x"626" => data <= "1000000000";
                when x"627" => data <= "1111110111";
                when x"628" => data <= "1000000000";
                when x"629" => data <= "1111110111";
                when x"62A" => data <= "1000000000";
                when x"62B" => data <= "1000000000";
                when x"62C" => data <= "1000000000";
                when x"62D" => data <= "1111110111";
                when x"62E" => data <= "1000000000";
                when x"62F" => data <= "1000000000";
                when x"630" => data <= "1000000000";
                when x"631" => data <= "1000000000";
                when x"632" => data <= "1111110111";
                when x"633" => data <= "1000000000";
                when x"634" => data <= "1000000000";
                when x"635" => data <= "1000000000";
                when x"636" => data <= "1111110111";
                when x"637" => data <= "1000000000";
                when x"638" => data <= "1111110111";
                when x"639" => data <= "1000000000";
                when x"63A" => data <= "1000000000";
                when x"63B" => data <= "0110000100";
                when x"63C" => data <= "1111110111";
                when x"63D" => data <= "1000000000";
                when x"63E" => data <= "1111110111";
                when x"63F" => data <= "1000000000";
                when x"640" => data <= "0101100101";
                when x"641" => data <= "1000000000";
                when x"642" => data <= "1000000000";
                when x"643" => data <= "1000000000";
                when x"644" => data <= "1000000000";
                when x"645" => data <= "0001110011";
                when x"646" => data <= "1000000000";
                when x"647" => data <= "1000000000";
                when x"648" => data <= "1000000000";
                when x"649" => data <= "1000000000";
                when x"64A" => data <= "1000000000";
                when x"64B" => data <= "1000000000";
                when x"64C" => data <= "1111110111";
                when x"64D" => data <= "1000000000";
                when x"64E" => data <= "0101010000";
                when x"64F" => data <= "1000000000";
                when x"650" => data <= "1000000000";
                when x"651" => data <= "1000000000";
                when x"652" => data <= "1000000000";
                when x"653" => data <= "1111110111";
                when x"654" => data <= "1000000000";
                when x"655" => data <= "1000000000";
                when x"656" => data <= "0101010000";
                when x"657" => data <= "1000000000";
                when x"658" => data <= "0101010000";
                when x"659" => data <= "1000110101";
                when x"65A" => data <= "1000000000";
                when x"65B" => data <= "1111110111";
                when x"65C" => data <= "1111110111";
                when x"65D" => data <= "1111110111";
                when x"65E" => data <= "1000000000";
                when x"65F" => data <= "0101010000";
                when x"660" => data <= "1111110111";
                when x"661" => data <= "0101010000";
                when x"662" => data <= "1000000000";
                when x"663" => data <= "1111110111";
                when x"664" => data <= "1000000000";
                when x"665" => data <= "1111110111";
                when x"666" => data <= "1111110111";
                when x"667" => data <= "1111110111";
                when x"668" => data <= "1111110111";
                when x"669" => data <= "1000000000";
                when x"66A" => data <= "1000000000";
                when x"66B" => data <= "1111110111";
                when x"66C" => data <= "1000000000";
                when x"66D" => data <= "1000000000";
                when x"66E" => data <= "1000000000";
                when x"66F" => data <= "1000000000";
                when x"670" => data <= "1000000000";
                when x"671" => data <= "1000000000";
                when x"672" => data <= "1111110111";
                when x"673" => data <= "1000000000";
                when x"674" => data <= "1000000000";
                when x"675" => data <= "0101100101";
                when x"676" => data <= "1000000000";
                when x"677" => data <= "0101100101";
                when x"678" => data <= "1111110111";
                when x"679" => data <= "1000000000";
                when x"67A" => data <= "1111110111";
                when x"67B" => data <= "1110101000";
                when x"67C" => data <= "1000000000";
                when x"67D" => data <= "1000000000";
                when x"67E" => data <= "1111110111";
                when x"67F" => data <= "1000000000";
                when x"680" => data <= "1111110111";
                when x"681" => data <= "1000000000";
                when x"682" => data <= "1000000000";
                when x"683" => data <= "1000000000";
                when x"684" => data <= "1000000000";
                when x"685" => data <= "1000000000";
                when x"686" => data <= "1111110111";
                when x"687" => data <= "1000000000";
                when x"688" => data <= "1111110111";
                when x"689" => data <= "1011010100";
                when x"68A" => data <= "1000000000";
                when x"68B" => data <= "1111110111";
                when x"68C" => data <= "1111110111";
                when x"68D" => data <= "0101010000";
                when x"68E" => data <= "1000000000";
                when x"68F" => data <= "1111110111";
                when x"690" => data <= "1000000000";
                when x"691" => data <= "1000000000";
                when x"692" => data <= "0010001000";
                when x"693" => data <= "0101111111";
                when x"694" => data <= "0101111111";
                when x"695" => data <= "1011111011";
                when x"696" => data <= "1111101101";
                when x"697" => data <= "0101111111";
                when x"698" => data <= "0100100000";
                when x"699" => data <= "1011111011";
                when x"69A" => data <= "0010001000";
                when x"69B" => data <= "0101111111";
                when x"69C" => data <= "1011111011";
                when x"69D" => data <= "0100010101";
                when x"69E" => data <= "0101111111";
                when x"69F" => data <= "0100010101";
                when x"6A0" => data <= "1111011000";
                when x"6A1" => data <= "0101001010";
                when x"6A2" => data <= "0010001000";
                when x"6A3" => data <= "1011111011";
                when x"6A4" => data <= "0010001000";
                when x"6A5" => data <= "0001101001";
                when x"6A6" => data <= "0010001000";
                when x"6A7" => data <= "1011111011";
                when x"6A8" => data <= "1111011000";
                when x"6A9" => data <= "0010001000";
                when x"6AA" => data <= "0010001000";
                when x"6AB" => data <= "0100010101";
                when x"6AC" => data <= "1111011000";
                when x"6AD" => data <= "1011111011";
                when x"6AE" => data <= "0010001000";
                when x"6AF" => data <= "1011111011";
                when x"6B0" => data <= "0010001000";
                when x"6B1" => data <= "1001110000";
                when x"6B2" => data <= "1011111011";
                when x"6B3" => data <= "1011111011";
                when x"6B4" => data <= "0100100000";
                when x"6B5" => data <= "0010001000";
                when x"6B6" => data <= "1011111011";
                when x"6B7" => data <= "0101111111";
                when x"6B8" => data <= "1111011000";
                when x"6B9" => data <= "0101111111";
                when x"6BA" => data <= "1011111011";
                when x"6BB" => data <= "0010001000";
                when x"6BC" => data <= "1011111011";
                when x"6BD" => data <= "1101010011";
                when x"6BE" => data <= "0000000011";
                when x"6BF" => data <= "1111011000";
                when x"6C0" => data <= "0010001000";
                when x"6C1" => data <= "0010001000";
                when x"6C2" => data <= "1011111011";
                when x"6C3" => data <= "1011111011";
                when x"6C4" => data <= "0010001000";
                when x"6C5" => data <= "1011111011";
                when x"6C6" => data <= "0101111111";
                when x"6C7" => data <= "0100100000";
                when x"6C8" => data <= "0101111111";
                when x"6C9" => data <= "1011111011";
                when x"6CA" => data <= "0010001000";
                when x"6CB" => data <= "1111011000";
                when x"6CC" => data <= "0101111111";
                when x"6CD" => data <= "0010001000";
                when x"6CE" => data <= "0101111111";
                when x"6CF" => data <= "1011111011";
                when x"6D0" => data <= "0100100000";
                when x"6D1" => data <= "0101111111";
                when x"6D2" => data <= "0101111111";
                when x"6D3" => data <= "1011001110";
                when x"6D4" => data <= "0101111111";
                when x"6D5" => data <= "0010001000";
                when x"6D6" => data <= "0110101011";
                when x"6D7" => data <= "1000101111";
                when x"6D8" => data <= "0101111111";
                when x"6D9" => data <= "1011111011";
                when x"6DA" => data <= "1011111011";
                when x"6DB" => data <= "0010001000";
                when x"6DC" => data <= "0101111111";
                when x"6DD" => data <= "1011111011";
                when x"6DE" => data <= "0010101010";
                when x"6DF" => data <= "0100110111";
                when x"6E0" => data <= "1001010010";
                when x"6E1" => data <= "1111111010";
                when x"6E2" => data <= "1111111010";
                when x"6E3" => data <= "0100000010";
                when x"6E4" => data <= "1010110011";
                when x"6E5" => data <= "0000100001";
                when x"6E6" => data <= "1111111010";
                when x"6E7" => data <= "0100000010";
                when x"6E8" => data <= "0011000000";
                when x"6E9" => data <= "1000111000";
                when x"6EA" => data <= "1001010010";
                when x"6EB" => data <= "0000100001";
                when x"6EC" => data <= "1001010010";
                when x"6ED" => data <= "0100000010";
                when x"6EE" => data <= "0110111100";
                when x"6EF" => data <= "1001010010";
                when x"6F0" => data <= "0000100001";
                when x"6F1" => data <= "0011000000";
                when x"6F2" => data <= "1111111010";
                when x"6F3" => data <= "1111111010";
                when x"6F4" => data <= "0010101010";
                when x"6F5" => data <= "0001001011";
                when x"6F6" => data <= "1011011001";
                when x"6F7" => data <= "0111010110";
                when x"6F8" => data <= "1001010010";
                when x"6F9" => data <= "1001010010";
                when x"6FA" => data <= "0111010110";
                when x"6FB" => data <= "0100110111";
                when x"6FC" => data <= "1000111000";
                when x"6FD" => data <= "0011000000";
                when x"6FE" => data <= "1000111000";
                when x"6FF" => data <= "1111001111";
                when x"700" => data <= "1111111010";
                when x"701" => data <= "0001001011";
                when x"702" => data <= "0100110111";
                when x"703" => data <= "0011000000";
                when x"704" => data <= "1111111010";
                when x"705" => data <= "1111111010";
                when x"706" => data <= "0101011101";
                when x"707" => data <= "1111111010";
                when x"708" => data <= "0000100001";
                when x"709" => data <= "1001010010";
                when x"70A" => data <= "1001010010";
                when x"70B" => data <= "1000001101";
                when x"70C" => data <= "0100000010";
                when x"70D" => data <= "0011000000";
                when x"70E" => data <= "0100000010";
                when x"70F" => data <= "1000111000";
                when x"710" => data <= "0111010110";
                when x"711" => data <= "0101011101";
                when x"712" => data <= "0011000000";
                when x"713" => data <= "0000100001";
                when x"714" => data <= "1111111010";
                when x"715" => data <= "0000100001";
                when x"716" => data <= "1111111010";
                when x"717" => data <= "0001111110";
                when x"718" => data <= "1111111010";
                when x"719" => data <= "1000001101";
                when x"71A" => data <= "1111111010";
                when x"71B" => data <= "0000010100";
                when x"71C" => data <= "1101110001";
                when x"71D" => data <= "1000111000";
                when x"71E" => data <= "0000100001";
                when x"71F" => data <= "1111111010";
                when x"720" => data <= "1000111000";
                when x"721" => data <= "0100000010";
                when x"722" => data <= "0100000010";
                when x"723" => data <= "1111111010";
                when x"724" => data <= "1001001000";
                when x"725" => data <= "0010000101";
                when x"726" => data <= "1110111111";
                when x"727" => data <= "1010101001";
                when x"728" => data <= "0000111011";
                when x"729" => data <= "0111001100";
                when x"72A" => data <= "0011101111";
                when x"72B" => data <= "0001100100";
                when x"72C" => data <= "0100101101";
                when x"72D" => data <= "1110111111";
                when x"72E" => data <= "0011011010";
                when x"72F" => data <= "1110111111";
                when x"730" => data <= "1110111111";
                when x"731" => data <= "1110111111";
                when x"732" => data <= "1110111111";
                when x"733" => data <= "1110111111";
                when x"734" => data <= "0100101101";
                when x"735" => data <= "1001111101";
                when x"736" => data <= "0010000101";
                when x"737" => data <= "0010000101";
                when x"738" => data <= "1101011110";
                when x"739" => data <= "1110111111";
                when x"73A" => data <= "1110111111";
                when x"73B" => data <= "1110111111";
                when x"73C" => data <= "1110111111";
                when x"73D" => data <= "1110111111";
                when x"73E" => data <= "1110111111";
                when x"73F" => data <= "1001111101";
                when x"740" => data <= "0100101101";
                when x"741" => data <= "1100110100";
                when x"742" => data <= "1110111111";
                when x"743" => data <= "1110111111";
                when x"744" => data <= "1110111111";
                when x"745" => data <= "1110111111";
                when x"746" => data <= "1001001000";
                when x"747" => data <= "1011110110";
                when x"748" => data <= "1001111101";
                when x"749" => data <= "1110111111";
                when x"74A" => data <= "0100101101";
                when x"74B" => data <= "1110111111";
                when x"74C" => data <= "1010101001";
                when x"74D" => data <= "1110111111";
                when x"74E" => data <= "1110111111";
                when x"74F" => data <= "0100101101";
                when x"750" => data <= "0011011010";
                when x"751" => data <= "1110111111";
                when x"752" => data <= "0011101111";
                when x"753" => data <= "1001001000";
                when x"754" => data <= "1011110110";
                when x"755" => data <= "1110111111";
                when x"756" => data <= "0010000000";
                when x"757" => data <= "0010000000";
                when x"758" => data <= "0101000010";
                when x"759" => data <= "1100110001";
                when x"75A" => data <= "0010000000";
                when x"75B" => data <= "1000010010";
                when x"75C" => data <= "0010000000";
                when x"75D" => data <= "1001111000";
                when x"75E" => data <= "0010000000";
                when x"75F" => data <= "1000100111";
                when x"760" => data <= "1011000110";
                when x"761" => data <= "0010000000";
                when x"762" => data <= "0101110111";
                when x"763" => data <= "0010000000";
                when x"764" => data <= "1000100111";
                when x"765" => data <= "0010000000";
                when x"766" => data <= "0010000000";
                when x"767" => data <= "0010000000";
                when x"768" => data <= "1100000100";
                when x"769" => data <= "1010101100";
                when x"76A" => data <= "0010000000";
                when x"76B" => data <= "0010000000";
                when x"76C" => data <= "0000001011";
                when x"76D" => data <= "1110111010";
                when x"76E" => data <= "0101110111";
                when x"76F" => data <= "0010000000";
                when x"770" => data <= "1111100101";
                when x"771" => data <= "1010101100";
                when x"772" => data <= "0010000000";
                when x"773" => data <= "0101110111";
                when x"774" => data <= "0101110111";
                when x"775" => data <= "0010000000";
                when x"776" => data <= "0101110111";
                when x"777" => data <= "0101000010";
                when x"778" => data <= "0101110111";
                when x"779" => data <= "1111010000";
                when x"77A" => data <= "1000010010";
                when x"77B" => data <= "1100110001";
                when x"77C" => data <= "0010000000";
                when x"77D" => data <= "0101110111";
                when x"77E" => data <= "0010000000";
                when x"77F" => data <= "0101000010";
                when x"780" => data <= "0101110111";
                when x"781" => data <= "1011110011";
                when x"782" => data <= "0010000000";
                when x"783" => data <= "1111010000";
                when x"784" => data <= "0010000000";
                when x"785" => data <= "0001010100";
                when x"786" => data <= "0010000000";
                when x"787" => data <= "0101110111";
                when x"788" => data <= "0010000000";
                when x"789" => data <= "0011101010";
                when x"78A" => data <= "1110111010";
                when x"78B" => data <= "0101000010";
                when x"78C" => data <= "0101110111";
                when x"78D" => data <= "0101000010";
                when x"78E" => data <= "0100101000";
                when x"78F" => data <= "0010000000";
                when x"790" => data <= "0010000000";
                when x"791" => data <= "0010000000";
                when x"792" => data <= "1100000100";
                when x"793" => data <= "0111111100";
                when x"794" => data <= "0010000000";
                when x"795" => data <= "0010000000";
                when x"796" => data <= "0010000000";
                when x"797" => data <= "0101110111";
                when x"798" => data <= "1000010010";
                when x"799" => data <= "0011011111";
                when x"79A" => data <= "0100101000";
                when x"79B" => data <= "0101000010";
                when x"79C" => data <= "1000010010";
                when x"79D" => data <= "0101110111";
                when x"79E" => data <= "1100000100";
                when x"79F" => data <= "0101000010";
                when x"7A0" => data <= "0010000000";
                when x"7A1" => data <= "1000100111";
                when x"7A2" => data <= "1111111111";
                when x"7A3" => data <= "1111111111";
                when x"7A4" => data <= "1111111111";
                when x"7A5" => data <= "1111111111";
                when x"7A6" => data <= "1111111111";
                when x"7A7" => data <= "1111111111";
                when x"7A8" => data <= "1111111111";
                when x"7A9" => data <= "1111111111";
                when x"7AA" => data <= "1111111111";
                when x"7AB" => data <= "1111111111";
                when x"7AC" => data <= "1111111111";
                when x"7AD" => data <= "1111111111";
                when x"7AE" => data <= "1111111111";
                when x"7AF" => data <= "1111111111";
                when x"7B0" => data <= "1111111111";
                when x"7B1" => data <= "1111111111";
                when x"7B2" => data <= "1111111111";
                when x"7B3" => data <= "1111111111";
                when x"7B4" => data <= "1111111111";
                when x"7B5" => data <= "1111111111";
                when x"7B6" => data <= "1111111111";
                when x"7B7" => data <= "1111111111";
                when x"7B8" => data <= "1111111111";
                when x"7B9" => data <= "1111111111";
                when x"7BA" => data <= "1111111111";
                when x"7BB" => data <= "1000001000";
                when x"7BC" => data <= "1111111111";
                when x"7BD" => data <= "1111111111";
                when x"7BE" => data <= "1111111111";
                when x"7BF" => data <= "1111111111";
                when x"7C0" => data <= "1111111111";
                when x"7C1" => data <= "1111111111";
                when x"7C2" => data <= "1111111111";
                when x"7C3" => data <= "1111111111";
                when x"7C4" => data <= "1111111111";
                when x"7C5" => data <= "1111111111";
                when x"7C6" => data <= "1111111111";
                when x"7C7" => data <= "1111111111";
                when x"7C8" => data <= "1111111111";
                when x"7C9" => data <= "1111111111";
                when x"7CA" => data <= "1111111111";
                when x"7CB" => data <= "1111111111";
                when x"7CC" => data <= "1111111111";
                when x"7CD" => data <= "1111111111";
                when x"7CE" => data <= "1111111111";
                when x"7CF" => data <= "1111111111";
                when x"7D0" => data <= "1111111111";
                when x"7D1" => data <= "1111111111";
                when x"7D2" => data <= "1111111111";
                when x"7D3" => data <= "1111111111";
                when x"7D4" => data <= "1111111111";
                when x"7D5" => data <= "1111111111";
                when x"7D6" => data <= "1111111111";
                when x"7D7" => data <= "1111111111";
                when x"7D8" => data <= "1111111111";
                when x"7D9" => data <= "1111111111";
                when x"7DA" => data <= "1111111111";
                when x"7DB" => data <= "1111111111";
                when x"7DC" => data <= "1111111111";
                when x"7DD" => data <= "1111111111";
                when x"7DE" => data <= "1111111111";
                when x"7DF" => data <= "1111111111";
                when x"7E0" => data <= "1111111111";
                when x"7E1" => data <= "1111111111";
                when x"7E2" => data <= "1111111111";
                when x"7E3" => data <= "1111111111";
                when x"7E4" => data <= "1111111111";
                when x"7E5" => data <= "1111111111";
                when x"7E6" => data <= "1111111111";
                when x"7E7" => data <= "1111111111";
                when x"7E8" => data <= "1111111111";
                when x"7E9" => data <= "1111111111";
                when x"7EA" => data <= "1111111111";
                when x"7EB" => data <= "1111111111";
                when x"7EC" => data <= "1111111111";
                when x"7ED" => data <= "1111111111";
                when x"7EE" => data <= "1111111111";
                when x"7EF" => data <= "1111111111";
                when x"7F0" => data <= "1111111111";
                when x"7F1" => data <= "1111111111";
                when x"7F2" => data <= "1111111111";
                when x"7F3" => data <= "1111111111";
                when x"7F4" => data <= "1111111111";
                when x"7F5" => data <= "1111111111";
                when x"7F6" => data <= "1111111111";
                when x"7F7" => data <= "1111111111";
                when x"7F8" => data <= "1111111111";
                when x"7F9" => data <= "1111111111";
                when x"7FA" => data <= "1111111111";
                when x"7FB" => data <= "1111111111";
                when x"7FC" => data <= "1111111111";
                when x"7FD" => data <= "1111111111";
                when x"7FE" => data <= "1111111111";
                when x"7FF" => data <= "1111111111";
                when x"800" => data <= "1111111111";
                when x"801" => data <= "1111111111";
                when x"802" => data <= "1111111111";
                when x"803" => data <= "1111111111";
                when x"804" => data <= "1111111111";
                when x"805" => data <= "1111111111";
                when x"806" => data <= "1111111111";
                when x"807" => data <= "1111111111";
                when x"808" => data <= "1111111111";
                when x"809" => data <= "1111111111";
                when x"80A" => data <= "1111111111";
                when x"80B" => data <= "1111111111";
                when x"80C" => data <= "1111111111";
                when x"80D" => data <= "1111111111";
                when x"80E" => data <= "1111111111";
                when x"80F" => data <= "1111111111";
                when x"810" => data <= "1111111111";
                when x"811" => data <= "1111111111";
                when x"812" => data <= "1111111111";
                when x"813" => data <= "1111111111";
                when x"814" => data <= "1111111111";
                when x"815" => data <= "1111111111";
                when x"816" => data <= "1111111111";
                when x"817" => data <= "1111111111";
                when x"818" => data <= "1111111111";
                when x"819" => data <= "1111111111";
                when x"81A" => data <= "1111111111";
                when x"81B" => data <= "1111111111";
                when x"81C" => data <= "1111111111";
                when x"81D" => data <= "1111111111";
                when x"81E" => data <= "1111111111";
                when x"81F" => data <= "1111111111";
                when x"820" => data <= "1111111111";
                when x"821" => data <= "1111111111";
                when x"822" => data <= "1111111111";
                when x"823" => data <= "1111111111";
                when x"824" => data <= "1111111111";
                when x"825" => data <= "1111111111";
                when x"826" => data <= "1111111111";
                when x"827" => data <= "1111111111";
                when x"828" => data <= "1111111111";
                when x"829" => data <= "1111111111";
                when x"82A" => data <= "1111111111";
                when x"82B" => data <= "1111111111";
                when x"82C" => data <= "1111111111";
                when x"82D" => data <= "1111111111";
                when x"82E" => data <= "1111111111";
                when x"82F" => data <= "1111111111";
                when x"830" => data <= "1111111111";
                when x"831" => data <= "1111111111";
                when x"832" => data <= "1111111111";
                when x"833" => data <= "1111111111";
                when x"834" => data <= "1111111111";
                when x"835" => data <= "1111111111";
                when x"836" => data <= "1111111111";
                when x"837" => data <= "1111111111";
                when x"838" => data <= "1111111111";
                when x"839" => data <= "1111111111";
                when x"83A" => data <= "1111111111";
                when x"83B" => data <= "1111111111";
                when x"83C" => data <= "1111111111";
                when x"83D" => data <= "1111111111";
                when x"83E" => data <= "1111111111";
                when x"83F" => data <= "1111111111";
                when x"840" => data <= "1111111111";
                when x"841" => data <= "1111111111";
                when x"842" => data <= "1111111111";
                when x"843" => data <= "1111111111";
                when x"844" => data <= "1111111111";
                when x"845" => data <= "1111111111";
                when x"846" => data <= "1111111111";
                when x"847" => data <= "1111111111";
                when x"848" => data <= "1111111111";
                when x"849" => data <= "1111111111";
                when x"84A" => data <= "1111111111";
                when x"84B" => data <= "1111111111";
                when x"84C" => data <= "1111111111";
                when x"84D" => data <= "1111111111";
                when x"84E" => data <= "1111111111";
                when x"84F" => data <= "1111111111";
                when x"850" => data <= "1111111111";
                when x"851" => data <= "1111111111";
                when x"852" => data <= "1111111111";
                when x"853" => data <= "1111111111";
                when x"854" => data <= "1111111111";
                when x"855" => data <= "1111111111";
                when x"856" => data <= "1111111111";
                when x"857" => data <= "1111111111";
                when x"858" => data <= "1111111111";
                when x"859" => data <= "1111111111";
                when x"85A" => data <= "1111111111";
                when x"85B" => data <= "1111111111";
                when x"85C" => data <= "1111111111";
                when x"85D" => data <= "1111111111";
                when x"85E" => data <= "1111111111";
                when x"85F" => data <= "1111111111";
                when x"860" => data <= "1111111111";
                when x"861" => data <= "1111111111";
                when x"862" => data <= "1111111111";
                when x"863" => data <= "1111111111";
                when x"864" => data <= "1111111111";
                when x"865" => data <= "1111111111";
                when x"866" => data <= "1111111111";
                when x"867" => data <= "1011101001";
                when x"868" => data <= "1111111111";
                when x"869" => data <= "1111111111";
                when x"86A" => data <= "1111111111";
                when x"86B" => data <= "1111111111";
                when x"86C" => data <= "1111111111";
                when x"86D" => data <= "1111111111";
                when x"86E" => data <= "1111111111";
                when x"86F" => data <= "1111111111";
                when x"870" => data <= "1111111111";
                when x"871" => data <= "1111111111";
                when x"872" => data <= "1111111111";
                when x"873" => data <= "1111111111";
                when x"874" => data <= "1111111111";
                when x"875" => data <= "1111111111";
                when x"876" => data <= "1111111111";
                when x"877" => data <= "1111111111";
                when x"878" => data <= "1111111111";
                when x"879" => data <= "1111111111";
                when x"87A" => data <= "1111111111";
                when x"87B" => data <= "1111111111";
                when x"87C" => data <= "1111111111";
                when x"87D" => data <= "1111111111";
                when x"87E" => data <= "1111111111";
                when x"87F" => data <= "1111111111";
                when x"880" => data <= "1111111111";
                when x"881" => data <= "1111111111";
                when x"882" => data <= "1111111111";
                when x"883" => data <= "1111111111";
                when x"884" => data <= "1111111111";
                when x"885" => data <= "1111111111";
                when x"886" => data <= "1111111111";
                when x"887" => data <= "1111111111";
                when x"888" => data <= "1111111111";
                when x"889" => data <= "1111111111";
                when x"88A" => data <= "1111111111";
                when x"88B" => data <= "1111111111";
                when x"88C" => data <= "1111111111";
                when x"88D" => data <= "1111111111";
                when x"88E" => data <= "1111111111";
                when x"88F" => data <= "1111111111";
                when x"890" => data <= "1111111111";
                when x"891" => data <= "1111111111";
                when x"892" => data <= "1111111111";
                when x"893" => data <= "1111111111";
                when x"894" => data <= "1111111111";
                when x"895" => data <= "1111111111";
                when x"896" => data <= "1111111111";
                when x"897" => data <= "1111111111";
                when x"898" => data <= "1111111111";
                when x"899" => data <= "1111111111";
                when x"89A" => data <= "1111111111";
                when x"89B" => data <= "1111111111";
                when x"89C" => data <= "1111111111";
                when x"89D" => data <= "1111111111";
                when x"89E" => data <= "1111111111";
                when x"89F" => data <= "1111111111";
                when x"8A0" => data <= "1111111111";
                when x"8A1" => data <= "1111111111";
                when x"8A2" => data <= "1111111111";
                when x"8A3" => data <= "1111111111";
                when x"8A4" => data <= "1111111111";
                when x"8A5" => data <= "1111111111";
                when x"8A6" => data <= "1111111111";
                when x"8A7" => data <= "1111111111";
                when x"8A8" => data <= "1111111111";
                when x"8A9" => data <= "1111111111";
                when x"8AA" => data <= "1111111111";
                when x"8AB" => data <= "1111111111";
                when x"8AC" => data <= "1111111111";
                when x"8AD" => data <= "1111111111";
                when x"8AE" => data <= "1111111111";
                when x"8AF" => data <= "1111111111";
                when x"8B0" => data <= "1111111111";
                when x"8B1" => data <= "1111111111";
                when x"8B2" => data <= "1111111111";
                when x"8B3" => data <= "1111111111";
                when x"8B4" => data <= "1111111111";
                when x"8B5" => data <= "1111111111";
                when x"8B6" => data <= "1111111111";
                when x"8B7" => data <= "1111111111";
                when x"8B8" => data <= "1111111111";
                when x"8B9" => data <= "1111111111";
                when x"8BA" => data <= "1111111111";
                when x"8BB" => data <= "1111111111";
                when x"8BC" => data <= "1111111111";
                when x"8BD" => data <= "1111111111";
                when x"8BE" => data <= "1111111111";
                when x"8BF" => data <= "1111111111";
                when x"8C0" => data <= "1111111111";
                when x"8C1" => data <= "1111111111";
                when x"8C2" => data <= "1111111111";
                when x"8C3" => data <= "1111111111";
                when x"8C4" => data <= "1111111111";
                when x"8C5" => data <= "1111111111";
                when x"8C6" => data <= "1111111111";
                when x"8C7" => data <= "1111111111";
                when x"8C8" => data <= "1111111111";
                when x"8C9" => data <= "1111111111";
                when x"8CA" => data <= "1111111111";
                when x"8CB" => data <= "1111111111";
                when x"8CC" => data <= "1111111111";
                when x"8CD" => data <= "1111111111";
                when x"8CE" => data <= "1111111111";
                when x"8CF" => data <= "1111111111";
                when x"8D0" => data <= "1111111111";
                when x"8D1" => data <= "1000001000";
                when x"8D2" => data <= "1111111111";
                when x"8D3" => data <= "1111111111";
                when x"8D4" => data <= "1111111111";
                when x"8D5" => data <= "1111111111";
                when x"8D6" => data <= "1111111111";
                when x"8D7" => data <= "1000001000";
                when x"8D8" => data <= "1111111111";
                when x"8D9" => data <= "1111111111";
                when x"8DA" => data <= "1111111111";
                when x"8DB" => data <= "1111111111";
                when x"8DC" => data <= "1111111111";
                when x"8DD" => data <= "1111111111";
                when x"8DE" => data <= "1111001010";
                when x"8DF" => data <= "1111111111";
                when x"8E0" => data <= "1111111111";
                when x"8E1" => data <= "1000001000";
                when x"8E2" => data <= "1111111111";
                when x"8E3" => data <= "1111111111";
                when x"8E4" => data <= "1111111111";
                when x"8E5" => data <= "1111111111";
                when x"8E6" => data <= "1111111111";
                when x"8E7" => data <= "1111111111";
                when x"8E8" => data <= "1111111111";
                when x"8E9" => data <= "1111111111";
                when x"8EA" => data <= "1111111111";
                when x"8EB" => data <= "1111111111";
                when x"8EC" => data <= "1111111111";
                when x"8ED" => data <= "1111111111";
                when x"8EE" => data <= "1111111111";
                when x"8EF" => data <= "1111111111";
                when x"8F0" => data <= "1111111111";
                when x"8F1" => data <= "1111111111";
                when x"8F2" => data <= "1111111111";
                when x"8F3" => data <= "1111111111";
                when x"8F4" => data <= "1111111111";
                when x"8F5" => data <= "1111111111";
                when x"8F6" => data <= "1111111111";
                when x"8F7" => data <= "1111111111";
                when x"8F8" => data <= "1111111111";
                when x"8F9" => data <= "1111111111";
                when x"8FA" => data <= "1111111111";
                when x"8FB" => data <= "1111111111";
                when x"8FC" => data <= "1111111111";
                when x"8FD" => data <= "1111111111";
                when x"8FE" => data <= "1111111111";
                when x"8FF" => data <= "1111111111";
                when x"900" => data <= "1111111111";
                when x"901" => data <= "1111111111";
                when x"902" => data <= "1111111111";
                when x"903" => data <= "1111111111";
                when x"904" => data <= "1111111111";
                when x"905" => data <= "1111111111";
                when x"906" => data <= "1111111111";
                when x"907" => data <= "1111111111";
                when x"908" => data <= "1111111111";
                when x"909" => data <= "1111111111";
                when x"90A" => data <= "1111111111";
                when x"90B" => data <= "1111111111";
                when x"90C" => data <= "1111111111";
                when x"90D" => data <= "1111111111";
                when x"90E" => data <= "1111111111";
                when x"90F" => data <= "1111111111";
                when x"910" => data <= "1111111111";
                when x"911" => data <= "1111111111";
                when x"912" => data <= "1111111111";
                when x"913" => data <= "1111111111";
                when x"914" => data <= "1111111111";
                when x"915" => data <= "1111111111";
                when x"916" => data <= "1111111111";
                when x"917" => data <= "1111111111";
                when x"918" => data <= "1111111111";
                when x"919" => data <= "1111111111";
                when x"91A" => data <= "1111111111";
                when x"91B" => data <= "1111111111";
                when x"91C" => data <= "1111111111";
                when x"91D" => data <= "1111111111";
                when x"91E" => data <= "1111111111";
                when x"91F" => data <= "1111111111";
                when x"920" => data <= "1111111111";
                when x"921" => data <= "1111111111";
                when x"922" => data <= "1111111111";
                when x"923" => data <= "1111111111";
                when x"924" => data <= "1111111111";
                when x"925" => data <= "1111111111";
                when x"926" => data <= "1111111111";
                when x"927" => data <= "1111111111";
                when x"928" => data <= "1111111111";
                when x"929" => data <= "1111111111";
                when x"92A" => data <= "1111111111";
                when x"92B" => data <= "1111111111";
                when x"92C" => data <= "1111111111";
                when x"92D" => data <= "1111111111";
                when x"92E" => data <= "1111111111";
                when x"92F" => data <= "1111111111";
                when x"930" => data <= "1111111111";
                when x"931" => data <= "1111111111";
                when x"932" => data <= "1111111111";
                when x"933" => data <= "1111111111";
                when x"934" => data <= "1111111111";
                when x"935" => data <= "1111111111";
                when x"936" => data <= "1111111111";
                when x"937" => data <= "1111111111";
                when x"938" => data <= "1111111111";
                when x"939" => data <= "1111111111";
                when x"93A" => data <= "1111111111";
                when x"93B" => data <= "1111111111";
                when x"93C" => data <= "1111111111";
                when x"93D" => data <= "1111111111";
                when x"93E" => data <= "1111111111";
                when x"93F" => data <= "1111111111";
                when x"940" => data <= "1111111111";
                when x"941" => data <= "1111111111";
                when x"942" => data <= "1111111111";
                when x"943" => data <= "1111111111";
                when x"944" => data <= "1111111111";
                when x"945" => data <= "1111111111";
                when x"946" => data <= "1111111111";
                when x"947" => data <= "1111111111";
                when x"948" => data <= "1111111111";
                when x"949" => data <= "1111111111";
                when x"94A" => data <= "1111111111";
                when x"94B" => data <= "1111111111";
                when x"94C" => data <= "1111111111";
                when x"94D" => data <= "1111111111";
                when x"94E" => data <= "1111111111";
                when x"94F" => data <= "1111111111";
                when x"950" => data <= "1111111111";
                when x"951" => data <= "1111111111";
                when x"952" => data <= "1111111111";
                when x"953" => data <= "1111111111";
                when x"954" => data <= "1111111111";
                when x"955" => data <= "1111111111";
                when x"956" => data <= "1111111111";
                when x"957" => data <= "1111111111";
                when x"958" => data <= "1111111111";
                when x"959" => data <= "1111111111";
                when x"95A" => data <= "1111111111";
                when x"95B" => data <= "1111111111";
                when x"95C" => data <= "1111111111";
                when x"95D" => data <= "1111111111";
                when x"95E" => data <= "1111111111";
                when x"95F" => data <= "1111111111";
                when x"960" => data <= "1111111111";
                when x"961" => data <= "1111111111";
                when x"962" => data <= "1111111111";
                when x"963" => data <= "1111111111";
                when x"964" => data <= "1111111111";
                when x"965" => data <= "1111111111";
                when x"966" => data <= "1111111111";
                when x"967" => data <= "1111111111";
                when x"968" => data <= "1111111111";
                when x"969" => data <= "1111111111";
                when x"96A" => data <= "1111111111";
                when x"96B" => data <= "1111111111";
                when x"96C" => data <= "1111111111";
                when x"96D" => data <= "1111111111";
                when x"96E" => data <= "1111111111";
                when x"96F" => data <= "1111111111";
                when x"970" => data <= "1111111111";
                when x"971" => data <= "1111111111";
                when x"972" => data <= "1111111111";
                when x"973" => data <= "1111111111";
                when x"974" => data <= "0010011010";
                when x"975" => data <= "1111111111";
                when x"976" => data <= "1111111111";
                when x"977" => data <= "1111111111";
                when x"978" => data <= "1111111111";
                when x"979" => data <= "1111111111";
                when x"97A" => data <= "1111111111";
                when x"97B" => data <= "1111111111";
                when x"97C" => data <= "1111111111";
                when x"97D" => data <= "1111111111";
                when x"97E" => data <= "1111111111";
                when x"97F" => data <= "1111111111";
                when x"980" => data <= "1111111111";
                when x"981" => data <= "1111111111";
                when x"982" => data <= "1111111111";
                when x"983" => data <= "1111111111";
                when x"984" => data <= "1111111111";
                when x"985" => data <= "1111111111";
                when x"986" => data <= "1111111111";
                when x"987" => data <= "1111111111";
                when x"988" => data <= "1111111111";
                when x"989" => data <= "1111111111";
                when x"98A" => data <= "1111111111";
                when x"98B" => data <= "1111111111";
                when x"98C" => data <= "1111111111";
                when x"98D" => data <= "1111111111";
                when x"98E" => data <= "1111111111";
                when x"98F" => data <= "1111111111";
                when x"990" => data <= "1111111111";
                when x"991" => data <= "1111111111";
                when x"992" => data <= "1111111111";
                when x"993" => data <= "1111111111";
                when x"994" => data <= "1111111111";
                when x"995" => data <= "1111111111";
                when x"996" => data <= "1111111111";
                when x"997" => data <= "1111111111";
                when x"998" => data <= "1111111111";
                when x"999" => data <= "1111111111";
                when x"99A" => data <= "1111111111";
                when x"99B" => data <= "1111111111";
                when x"99C" => data <= "1111111111";
                when x"99D" => data <= "1111111111";
                when x"99E" => data <= "1111111111";
                when x"99F" => data <= "1111111111";
                when x"9A0" => data <= "1111111111";
                when x"9A1" => data <= "1111111111";
                when x"9A2" => data <= "1111111111";
                when x"9A3" => data <= "1111111111";
                when x"9A4" => data <= "1111111111";
                when x"9A5" => data <= "1111111111";
                when x"9A6" => data <= "1111111111";
                when x"9A7" => data <= "1111111111";
                when x"9A8" => data <= "1111111111";
                when x"9A9" => data <= "1111111111";
                when x"9AA" => data <= "1111111111";
                when x"9AB" => data <= "1111111111";
                when x"9AC" => data <= "1111111111";
                when x"9AD" => data <= "1111111111";
                when x"9AE" => data <= "1111111111";
                when x"9AF" => data <= "1111111111";
                when x"9B0" => data <= "1111111111";
                when x"9B1" => data <= "1111111111";
                when x"9B2" => data <= "1111111111";
                when x"9B3" => data <= "1111111111";
                when x"9B4" => data <= "1111111111";
                when x"9B5" => data <= "1111111111";
                when x"9B6" => data <= "1111111111";
                when x"9B7" => data <= "1111111111";
                when x"9B8" => data <= "1111111111";
                when x"9B9" => data <= "1111111111";
                when x"9BA" => data <= "1111111111";
                when x"9BB" => data <= "1111111111";
                when x"9BC" => data <= "1111111111";
                when x"9BD" => data <= "1111111111";
                when x"9BE" => data <= "1111111111";
                when x"9BF" => data <= "1111111111";
                when x"9C0" => data <= "1111111111";
                when x"9C1" => data <= "1111111111";
                when x"9C2" => data <= "1111111111";
                when x"9C3" => data <= "1111111111";
                when x"9C4" => data <= "1111111111";
                when x"9C5" => data <= "1111111111";
                when x"9C6" => data <= "1111111111";
                when x"9C7" => data <= "1111111111";
                when x"9C8" => data <= "1111111111";
                when x"9C9" => data <= "1111111111";
                when x"9CA" => data <= "1111111111";
                when x"9CB" => data <= "1111111111";
                when x"9CC" => data <= "1111111111";
                when x"9CD" => data <= "1111111111";
                when x"9CE" => data <= "1111111111";
                when x"9CF" => data <= "1111111111";
                when x"9D0" => data <= "1111111111";
                when x"9D1" => data <= "1111111111";
                when x"9D2" => data <= "1111111111";
                when x"9D3" => data <= "1111111111";
                when x"9D4" => data <= "1111111111";
                when x"9D5" => data <= "1111111111";
                when x"9D6" => data <= "1111111111";
                when x"9D7" => data <= "1111111111";
                when x"9D8" => data <= "1111111111";
                when x"9D9" => data <= "1111111111";
                when x"9DA" => data <= "1111111111";
                when x"9DB" => data <= "1111111111";
                when x"9DC" => data <= "1111111111";
                when x"9DD" => data <= "1111111111";
                when x"9DE" => data <= "1111111111";
                when x"9DF" => data <= "1111111111";
                when x"9E0" => data <= "1111111111";
                when x"9E1" => data <= "1111111111";
                when x"9E2" => data <= "1111111111";
                when x"9E3" => data <= "1111111111";
                when x"9E4" => data <= "1111111111";
                when x"9E5" => data <= "1111111111";
                when x"9E6" => data <= "1111111111";
                when x"9E7" => data <= "1111111111";
                when x"9E8" => data <= "1111111111";
                when x"9E9" => data <= "1111111111";
                when x"9EA" => data <= "1111111111";
                when x"9EB" => data <= "1111111111";
                when x"9EC" => data <= "1111111111";
                when x"9ED" => data <= "1111111111";
                when x"9EE" => data <= "1111111111";
                when x"9EF" => data <= "1111111111";
                when x"9F0" => data <= "1111111111";
                when x"9F1" => data <= "1111111111";
                when x"9F2" => data <= "1111111111";
                when x"9F3" => data <= "1111111111";
                when x"9F4" => data <= "1111111111";
                when x"9F5" => data <= "1111111111";
                when x"9F6" => data <= "1111111111";
                when x"9F7" => data <= "1111111111";
                when x"9F8" => data <= "1111111111";
                when x"9F9" => data <= "1111111111";
                when x"9FA" => data <= "1111111111";
                when x"9FB" => data <= "1111111111";
                when x"9FC" => data <= "1111111111";
                when x"9FD" => data <= "1111111111";
                when x"9FE" => data <= "1111111111";
                when x"9FF" => data <= "1111111111";
                when x"A00" => data <= "1111111111";
                when x"A01" => data <= "1111111111";
                when x"A02" => data <= "1111111111";
                when x"A03" => data <= "1111111111";
                when x"A04" => data <= "1111111111";
                when x"A05" => data <= "1111111111";
                when x"A06" => data <= "1111111111";
                when x"A07" => data <= "1111111111";
                when x"A08" => data <= "1111111111";
                when x"A09" => data <= "1111111111";
                when x"A0A" => data <= "1111111111";
                when x"A0B" => data <= "1111111111";
                when x"A0C" => data <= "1111111111";
                when x"A0D" => data <= "1111111111";
                when x"A0E" => data <= "1111111111";
                when x"A0F" => data <= "1111111111";
                when x"A10" => data <= "1111111111";
                when x"A11" => data <= "1111111111";
                when x"A12" => data <= "1111111111";
                when x"A13" => data <= "1111111111";
                when x"A14" => data <= "1111111111";
                when x"A15" => data <= "1111111111";
                when x"A16" => data <= "1111111111";
                when x"A17" => data <= "1111111111";
                when x"A18" => data <= "1111111111";
                when x"A19" => data <= "1111111111";
                when x"A1A" => data <= "1111111111";
                when x"A1B" => data <= "1111111111";
                when x"A1C" => data <= "1111111111";
                when x"A1D" => data <= "1111111111";
                when x"A1E" => data <= "1111111111";
                when x"A1F" => data <= "1111111111";
                when x"A20" => data <= "1111111111";
                when x"A21" => data <= "1111111111";
                when x"A22" => data <= "1111111111";
                when x"A23" => data <= "1111111111";
                when x"A24" => data <= "1111111111";
                when x"A25" => data <= "1111111111";
                when x"A26" => data <= "1111111111";
                when x"A27" => data <= "1111111111";
                when x"A28" => data <= "1111111111";
                when x"A29" => data <= "1111111111";
                when x"A2A" => data <= "1111111111";
                when x"A2B" => data <= "1111111111";
                when x"A2C" => data <= "1111111111";
                when x"A2D" => data <= "1111111111";
                when x"A2E" => data <= "1111111111";
                when x"A2F" => data <= "1111111111";
                when x"A30" => data <= "1111111111";
                when x"A31" => data <= "1111111111";
                when x"A32" => data <= "1111111111";
                when x"A33" => data <= "1111111111";
                when x"A34" => data <= "1111111111";
                when x"A35" => data <= "1111111111";
                when x"A36" => data <= "1111111111";
                when x"A37" => data <= "1111111111";
                when x"A38" => data <= "1111111111";
                when x"A39" => data <= "1111111111";
                when x"A3A" => data <= "1111111111";
                when x"A3B" => data <= "1111111111";
                when x"A3C" => data <= "1111111111";
                when x"A3D" => data <= "1111111111";
                when x"A3E" => data <= "1111111111";
                when x"A3F" => data <= "1111111111";
                when x"A40" => data <= "1111111111";
                when x"A41" => data <= "1111111111";
                when x"A42" => data <= "1111111111";
                when x"A43" => data <= "1111111111";
                when x"A44" => data <= "1111111111";
                when x"A45" => data <= "1111111111";
                when x"A46" => data <= "1111111111";
                when x"A47" => data <= "1111111111";
                when x"A48" => data <= "1111111111";
                when x"A49" => data <= "1111111111";
                when x"A4A" => data <= "1111111111";
                when x"A4B" => data <= "1111111111";
                when x"A4C" => data <= "1111111111";
                when x"A4D" => data <= "1111111111";
                when x"A4E" => data <= "1111111111";
                when x"A4F" => data <= "1111111111";
                when x"A50" => data <= "1111111111";
                when x"A51" => data <= "1111111111";
                when x"A52" => data <= "1111111111";
                when x"A53" => data <= "1111111111";
                when x"A54" => data <= "1111111111";
                when x"A55" => data <= "1111111111";
                when x"A56" => data <= "1111111111";
                when x"A57" => data <= "1111111111";
                when x"A58" => data <= "1111111111";
                when x"A59" => data <= "1111111111";
                when x"A5A" => data <= "1111111111";
                when x"A5B" => data <= "1111111111";
                when x"A5C" => data <= "1111111111";
                when x"A5D" => data <= "1111111111";
                when x"A5E" => data <= "1111111111";
                when x"A5F" => data <= "1111111111";
                when x"A60" => data <= "1111111111";
                when x"A61" => data <= "1111111111";
                when x"A62" => data <= "1111111111";
                when x"A63" => data <= "1111111111";
                when x"A64" => data <= "1111111111";
                when x"A65" => data <= "1111111111";
                when x"A66" => data <= "1111111111";
                when x"A67" => data <= "1111111111";
                when x"A68" => data <= "1111111111";
                when x"A69" => data <= "1111111111";
                when x"A6A" => data <= "1111111111";
                when x"A6B" => data <= "1111111111";
                when x"A6C" => data <= "1111111111";
                when x"A6D" => data <= "1111111111";
                when x"A6E" => data <= "1111111111";
                when x"A6F" => data <= "1111111111";
                when x"A70" => data <= "1111111111";
                when x"A71" => data <= "1111111111";
                when x"A72" => data <= "1111111111";
                when x"A73" => data <= "1111111111";
                when x"A74" => data <= "1111111111";
                when x"A75" => data <= "1111111111";
                when x"A76" => data <= "1111111111";
                when x"A77" => data <= "1111111111";
                when x"A78" => data <= "1111111111";
                when x"A79" => data <= "1111111111";
                when x"A7A" => data <= "1111111111";
                when x"A7B" => data <= "1111111111";
                when x"A7C" => data <= "1111111111";
                when x"A7D" => data <= "1111111111";
                when x"A7E" => data <= "1111111111";
                when x"A7F" => data <= "1111111111";
                when x"A80" => data <= "1111111111";
                when x"A81" => data <= "1111111111";
                when x"A82" => data <= "1111111111";
                when x"A83" => data <= "1111111111";
                when x"A84" => data <= "1111111111";
                when x"A85" => data <= "1111111111";
                when x"A86" => data <= "1111111111";
                when x"A87" => data <= "1111111111";
                when x"A88" => data <= "1111111111";
                when x"A89" => data <= "0111010011";
                when x"A8A" => data <= "1111111111";
                when x"A8B" => data <= "1111111111";
                when x"A8C" => data <= "1000001000";
                when x"A8D" => data <= "1111111111";
                when x"A8E" => data <= "1111111111";
                when x"A8F" => data <= "1111111111";
                when x"A90" => data <= "1111111111";
                when x"A91" => data <= "1111111111";
                when x"A92" => data <= "1111111111";
                when x"A93" => data <= "1111111111";
                when x"A94" => data <= "1111111111";
                when x"A95" => data <= "1111111111";
                when x"A96" => data <= "1111111111";
                when x"A97" => data <= "1111111111";
                when x"A98" => data <= "1111111111";
                when x"A99" => data <= "1111111111";
                when x"A9A" => data <= "1111111111";
                when x"A9B" => data <= "1111111111";
                when x"A9C" => data <= "1111111111";
                when x"A9D" => data <= "1111111111";
                when x"A9E" => data <= "1111111111";
                when x"A9F" => data <= "1111111111";
                when x"AA0" => data <= "1111111111";
                when x"AA1" => data <= "1111111111";
                when x"AA2" => data <= "1111111111";
                when x"AA3" => data <= "1111111111";
                when x"AA4" => data <= "1111111111";
                when x"AA5" => data <= "1111111111";
                when x"AA6" => data <= "1111111111";
                when x"AA7" => data <= "1111111111";
                when x"AA8" => data <= "1111111111";
                when x"AA9" => data <= "1111111111";
                when x"AAA" => data <= "1111111111";
                when x"AAB" => data <= "1111111111";
                when x"AAC" => data <= "1111111111";
                when x"AAD" => data <= "1111111111";
                when x"AAE" => data <= "1111111111";
                when x"AAF" => data <= "1111111111";
                when x"AB0" => data <= "1111111111";
                when x"AB1" => data <= "1111111111";
                when x"AB2" => data <= "1111111111";
                when x"AB3" => data <= "1111111111";
                when x"AB4" => data <= "1111111111";
                when x"AB5" => data <= "1111111111";
                when x"AB6" => data <= "1111111111";
                when x"AB7" => data <= "1111111111";
                when x"AB8" => data <= "1111111111";
                when x"AB9" => data <= "1111111111";
                when x"ABA" => data <= "1111111111";
                when x"ABB" => data <= "1111111111";
                when x"ABC" => data <= "1111111111";
                when x"ABD" => data <= "1111111111";
                when x"ABE" => data <= "1111111111";
                when x"ABF" => data <= "1111111111";
                when x"AC0" => data <= "1111111111";
                when x"AC1" => data <= "1111001010";
                when x"AC2" => data <= "1111111111";
                when x"AC3" => data <= "1111111111";
                when x"AC4" => data <= "1111111111";
                when x"AC5" => data <= "1111111111";
                when x"AC6" => data <= "1111111111";
                when x"AC7" => data <= "1111111111";
                when x"AC8" => data <= "1111111111";
                when x"AC9" => data <= "1111111111";
                when x"ACA" => data <= "1111111111";
                when x"ACB" => data <= "1111111111";
                when x"ACC" => data <= "1111111111";
                when x"ACD" => data <= "1111111111";
                when x"ACE" => data <= "1111111111";
                when x"ACF" => data <= "1111111111";
                when x"AD0" => data <= "1111111111";
                when x"AD1" => data <= "1111111111";
                when x"AD2" => data <= "1111111111";
                when x"AD3" => data <= "1111111111";
                when x"AD4" => data <= "1111111111";
                when x"AD5" => data <= "1111111111";
                when x"AD6" => data <= "1111111111";
                when x"AD7" => data <= "1111111111";
                when x"AD8" => data <= "1111111111";
                when x"AD9" => data <= "1111111111";
                when x"ADA" => data <= "1111111111";
                when x"ADB" => data <= "1111111111";
                when x"ADC" => data <= "1111111111";
                when x"ADD" => data <= "1111111111";
                when x"ADE" => data <= "1111111111";
                when x"ADF" => data <= "1111111111";
                when x"AE0" => data <= "1111111111";
                when x"AE1" => data <= "1111111111";
                when x"AE2" => data <= "1111111111";
                when x"AE3" => data <= "1111111111";
                when x"AE4" => data <= "1111111111";
                when x"AE5" => data <= "1111111111";
                when x"AE6" => data <= "1111111111";
                when x"AE7" => data <= "1111111111";
                when x"AE8" => data <= "1111111111";
                when x"AE9" => data <= "1111111111";
                when x"AEA" => data <= "1111111111";
                when x"AEB" => data <= "1111111111";
                when x"AEC" => data <= "1111111111";
                when x"AED" => data <= "1111111111";
                when x"AEE" => data <= "1111111111";
                when x"AEF" => data <= "1111111111";
                when x"AF0" => data <= "0010101111";
                when x"AF1" => data <= "1111111111";
                when x"AF2" => data <= "1111111111";
                when x"AF3" => data <= "1111111111";
                when x"AF4" => data <= "1111111111";
                when x"AF5" => data <= "1111111111";
                when x"AF6" => data <= "1111111111";
                when x"AF7" => data <= "1111111111";
                when x"AF8" => data <= "1111111111";
                when x"AF9" => data <= "1111111111";
                when x"AFA" => data <= "1111111111";
                when x"AFB" => data <= "1111111111";
                when x"AFC" => data <= "1111111111";
                when x"AFD" => data <= "1111111111";
                when x"AFE" => data <= "1111111111";
                when x"AFF" => data <= "1111111111";
                when x"B00" => data <= "1111111111";
                when x"B01" => data <= "1111111111";
                when x"B02" => data <= "1111111111";
                when x"B03" => data <= "1111111111";
                when x"B04" => data <= "1111111111";
                when x"B05" => data <= "1111111111";
                when x"B06" => data <= "1111111111";
                when x"B07" => data <= "1111111111";
                when x"B08" => data <= "1111111111";
                when x"B09" => data <= "1111111111";
                when x"B0A" => data <= "1111111111";
                when x"B0B" => data <= "1111111111";
                when x"B0C" => data <= "1111111111";
                when x"B0D" => data <= "1111111111";
                when x"B0E" => data <= "1111111111";
                when x"B0F" => data <= "1111111111";
                when x"B10" => data <= "1111111111";
                when x"B11" => data <= "1111111111";
                when x"B12" => data <= "1111111111";
                when x"B13" => data <= "1111111111";
                when x"B14" => data <= "1111111111";
                when x"B15" => data <= "1111111111";
                when x"B16" => data <= "1111111111";
                when x"B17" => data <= "1111111111";
                when x"B18" => data <= "1111111111";
                when x"B19" => data <= "1111111111";
                when x"B1A" => data <= "1000001000";
                when x"B1B" => data <= "1111111111";
                when x"B1C" => data <= "1111111111";
                when x"B1D" => data <= "1111111111";
                when x"B1E" => data <= "1111111111";
                when x"B1F" => data <= "1111111111";
                when x"B20" => data <= "1111111111";
                when x"B21" => data <= "1111111111";
                when x"B22" => data <= "1111111111";
                when x"B23" => data <= "1111111111";
                when x"B24" => data <= "1111111111";
                when x"B25" => data <= "1111111111";
                when x"B26" => data <= "1111111111";
                when x"B27" => data <= "1111111111";
                when x"B28" => data <= "1111111111";
                when x"B29" => data <= "1111111111";
                when x"B2A" => data <= "1111111111";
                when x"B2B" => data <= "0001111011";
                when x"B2C" => data <= "1111111111";
                when x"B2D" => data <= "1111111111";
                when x"B2E" => data <= "1111111111";
                when x"B2F" => data <= "1111111111";
                when x"B30" => data <= "1111111111";
                when x"B31" => data <= "1111111111";
                when x"B32" => data <= "1111111111";
                when x"B33" => data <= "1111111111";
                when x"B34" => data <= "1111111111";
                when x"B35" => data <= "1111111111";
                when x"B36" => data <= "1111111111";
                when x"B37" => data <= "1111111111";
                when x"B38" => data <= "1111111111";
                when x"B39" => data <= "1111111111";
                when x"B3A" => data <= "1111111111";
                when x"B3B" => data <= "1111111111";
                when x"B3C" => data <= "1111111111";
                when x"B3D" => data <= "1111111111";
                when x"B3E" => data <= "1111111111";
                when x"B3F" => data <= "1111111111";
                when x"B40" => data <= "1111111111";
                when x"B41" => data <= "1111111111";
                when x"B42" => data <= "1111111111";
                when x"B43" => data <= "1111111111";
                when x"B44" => data <= "1111111111";
                when x"B45" => data <= "1111111111";
                when x"B46" => data <= "1111111111";
                when x"B47" => data <= "1111111111";
                when x"B48" => data <= "1111111111";
                when x"B49" => data <= "1111111111";
                when x"B4A" => data <= "1111111111";
                when x"B4B" => data <= "1111111111";
                when x"B4C" => data <= "1111111111";
                when x"B4D" => data <= "1111111111";
                when x"B4E" => data <= "1111111111";
                when x"B4F" => data <= "1111111111";
                when x"B50" => data <= "1111111111";
                when x"B51" => data <= "1111111111";
                when x"B52" => data <= "1111111111";
                when x"B53" => data <= "1111111111";
                when x"B54" => data <= "1111111111";
                when x"B55" => data <= "1111111111";
                when x"B56" => data <= "1111111111";
                when x"B57" => data <= "1111111111";
                when x"B58" => data <= "1111111111";
                when x"B59" => data <= "1111111111";
                when x"B5A" => data <= "1111111111";
                when x"B5B" => data <= "1111111111";
                when x"B5C" => data <= "1111111111";
                when x"B5D" => data <= "1111111111";
                when x"B5E" => data <= "1111111111";
                when x"B5F" => data <= "1111111111";
                when x"B60" => data <= "1111111111";
                when x"B61" => data <= "1111111111";
                when x"B62" => data <= "1111111111";
                when x"B63" => data <= "1111111111";
                when x"B64" => data <= "1111111111";
                when x"B65" => data <= "1111111111";
                when x"B66" => data <= "1111111111";
                when x"B67" => data <= "1111111111";
                when x"B68" => data <= "1111111111";
                when x"B69" => data <= "1111111111";
                when x"B6A" => data <= "1111111111";
                when x"B6B" => data <= "1111111111";
                when x"B6C" => data <= "1111111111";
                when x"B6D" => data <= "1111111111";
                when x"B6E" => data <= "1111111111";
                when x"B6F" => data <= "1111111111";
                when x"B70" => data <= "1111111111";
                when x"B71" => data <= "1111111111";
                when x"B72" => data <= "1111111111";
                when x"B73" => data <= "1111111111";
                when x"B74" => data <= "1111111111";
                when x"B75" => data <= "1111111111";
                when x"B76" => data <= "1111111111";
                when x"B77" => data <= "1111111111";
                when x"B78" => data <= "1111111111";
                when x"B79" => data <= "1111111111";
                when x"B7A" => data <= "1111111111";
                when x"B7B" => data <= "1111111111";
                when x"B7C" => data <= "1111111111";
                when x"B7D" => data <= "1111111111";
                when x"B7E" => data <= "1111111111";
                when x"B7F" => data <= "1111111111";
                when x"B80" => data <= "1111111111";
                when x"B81" => data <= "1111111111";
                when x"B82" => data <= "1111111111";
                when x"B83" => data <= "1111111111";
                when x"B84" => data <= "1111111111";
                when x"B85" => data <= "1111111111";
                when x"B86" => data <= "1111111111";
                when x"B87" => data <= "1111111111";
                when x"B88" => data <= "1111111111";
                when x"B89" => data <= "1111111111";
                when x"B8A" => data <= "1111111111";
                when x"B8B" => data <= "1111111111";
                when x"B8C" => data <= "1111111111";
                when x"B8D" => data <= "1111111111";
                when x"B8E" => data <= "1111111111";
                when x"B8F" => data <= "1111111111";
                when x"B90" => data <= "1111111111";
                when x"B91" => data <= "1111111111";
                when x"B92" => data <= "1111111111";
                when x"B93" => data <= "1111111111";
                when x"B94" => data <= "1111111111";
                when x"B95" => data <= "1111111111";
                when x"B96" => data <= "1111111111";
                when x"B97" => data <= "1111111111";
                when x"B98" => data <= "1111111111";
                when x"B99" => data <= "1111111111";
                when x"B9A" => data <= "1111111111";
                when x"B9B" => data <= "1111111111";
                when x"B9C" => data <= "1111111111";
                when x"B9D" => data <= "1111111111";
                when x"B9E" => data <= "1111111111";
                when x"B9F" => data <= "1111111111";
                when x"BA0" => data <= "1111111111";
                when x"BA1" => data <= "1111111111";
                when x"BA2" => data <= "1111111111";
                when x"BA3" => data <= "1111111111";
                when x"BA4" => data <= "1111111111";
                when x"BA5" => data <= "1111111111";
                when x"BA6" => data <= "1111111111";
                when x"BA7" => data <= "1111111111";
                when x"BA8" => data <= "1111111111";
                when x"BA9" => data <= "1111111111";
                when x"BAA" => data <= "1111111111";
                when x"BAB" => data <= "1111111111";
                when x"BAC" => data <= "1111111111";
                when x"BAD" => data <= "1111111111";
                when x"BAE" => data <= "1111111111";
                when x"BAF" => data <= "1111111111";
                when x"BB0" => data <= "1111111111";
                when x"BB1" => data <= "1111111111";
                when x"BB2" => data <= "1111111111";
                when x"BB3" => data <= "1111111111";
                when x"BB4" => data <= "1111111111";
                when x"BB5" => data <= "1111111111";
                when x"BB6" => data <= "1111111111";
                when x"BB7" => data <= "1111111111";
                when x"BB8" => data <= "1111111111";
                when x"BB9" => data <= "1111111111";
                when x"BBA" => data <= "1111111111";
                when x"BBB" => data <= "1111111111";
                when x"BBC" => data <= "1111111111";
                when x"BBD" => data <= "1111111111";
                when x"BBE" => data <= "1111111111";
                when x"BBF" => data <= "1111111111";
                when x"BC0" => data <= "1111111111";
                when x"BC1" => data <= "1111111111";
                when x"BC2" => data <= "1111111111";
                when x"BC3" => data <= "1111111111";
                when x"BC4" => data <= "1111111111";
                when x"BC5" => data <= "1111111111";
                when x"BC6" => data <= "1111111111";
                when x"BC7" => data <= "1111111111";
                when x"BC8" => data <= "1111111111";
                when x"BC9" => data <= "1111111111";
                when x"BCA" => data <= "1111111111";
                when x"BCB" => data <= "1111111111";
                when x"BCC" => data <= "1111111111";
                when x"BCD" => data <= "1111111111";
                when x"BCE" => data <= "1111111111";
                when x"BCF" => data <= "1111111111";
                when x"BD0" => data <= "1111111111";
                when x"BD1" => data <= "1111111111";
                when x"BD2" => data <= "1111111111";
                when x"BD3" => data <= "1111111111";
                when x"BD4" => data <= "1111111111";
                when x"BD5" => data <= "1111111111";
                when x"BD6" => data <= "1111111111";
                when x"BD7" => data <= "1111111111";
                when x"BD8" => data <= "1111111111";
                when x"BD9" => data <= "1111111111";
                when x"BDA" => data <= "1111111111";
                when x"BDB" => data <= "1111111111";
                when x"BDC" => data <= "1111111111";
                when x"BDD" => data <= "1111111111";
                when x"BDE" => data <= "1111111111";
                when x"BDF" => data <= "1111111111";
                when x"BE0" => data <= "1111111111";
                when x"BE1" => data <= "1111111111";
                when x"BE2" => data <= "1111111111";
                when x"BE3" => data <= "1111111111";
                when x"BE4" => data <= "1111111111";
                when x"BE5" => data <= "1111111111";
                when x"BE6" => data <= "1111111111";
                when x"BE7" => data <= "1111111111";
                when x"BE8" => data <= "1111111111";
                when x"BE9" => data <= "1111111111";
                when x"BEA" => data <= "1111111111";
                when x"BEB" => data <= "1111111111";
                when x"BEC" => data <= "1001010111";
                when x"BED" => data <= "1111111111";
                when x"BEE" => data <= "1111111111";
                when x"BEF" => data <= "1111111111";
                when x"BF0" => data <= "1111111111";
                when x"BF1" => data <= "1111111111";
                when x"BF2" => data <= "1111111111";
                when x"BF3" => data <= "1111111111";
                when x"BF4" => data <= "1111111111";
                when x"BF5" => data <= "1111111111";
                when x"BF6" => data <= "1111111111";
                when x"BF7" => data <= "1111111111";
                when x"BF8" => data <= "1111111111";
                when x"BF9" => data <= "1111111111";
                when x"BFA" => data <= "1111111111";
                when x"BFB" => data <= "1111111111";
                when x"BFC" => data <= "1111111111";
                when x"BFD" => data <= "1111111111";
                when x"BFE" => data <= "1111111111";
                when x"BFF" => data <= "1111111111";
                when x"C00" => data <= "1111111111";
                when x"C01" => data <= "1111111111";
                when x"C02" => data <= "1111111111";
                when x"C03" => data <= "1111111111";
                when x"C04" => data <= "1111111111";
                when x"C05" => data <= "1111111111";
                when x"C06" => data <= "1111111111";
                when x"C07" => data <= "1111111111";
                when x"C08" => data <= "1111111111";
                when x"C09" => data <= "1111111111";
                when x"C0A" => data <= "1111111111";
                when x"C0B" => data <= "1111111111";
                when x"C0C" => data <= "1111111111";
                when x"C0D" => data <= "1111111111";
                when x"C0E" => data <= "1111111111";
                when x"C0F" => data <= "1111111111";
                when x"C10" => data <= "1111111111";
                when x"C11" => data <= "1111111111";
                when x"C12" => data <= "1111111111";
                when x"C13" => data <= "1111111111";
                when x"C14" => data <= "1111111111";
                when x"C15" => data <= "1111111111";
                when x"C16" => data <= "1111111111";
                when x"C17" => data <= "1111111111";
                when x"C18" => data <= "1111111111";
                when x"C19" => data <= "1111111111";
                when x"C1A" => data <= "1111111111";
                when x"C1B" => data <= "1111111111";
                when x"C1C" => data <= "1111111111";
                when x"C1D" => data <= "1111111111";
                when x"C1E" => data <= "1111111111";
                when x"C1F" => data <= "1111111111";
                when x"C20" => data <= "1111111111";
                when x"C21" => data <= "1111111111";
                when x"C22" => data <= "1111111111";
                when x"C23" => data <= "1111111111";
                when x"C24" => data <= "1111111111";
                when x"C25" => data <= "1111111111";
                when x"C26" => data <= "1111111111";
                when x"C27" => data <= "1111111111";
                when x"C28" => data <= "1111111111";
                when x"C29" => data <= "1111111111";
                when x"C2A" => data <= "0100000111";
                when x"C2B" => data <= "1111111111";
                when x"C2C" => data <= "1111111111";
                when x"C2D" => data <= "1111111111";
                when x"C2E" => data <= "1111111111";
                when x"C2F" => data <= "1111111111";
                when x"C30" => data <= "1111111111";
                when x"C31" => data <= "1111111111";
                when x"C32" => data <= "1111111111";
                when x"C33" => data <= "1111111111";
                when x"C34" => data <= "1111111111";
                when x"C35" => data <= "1111111111";
                when x"C36" => data <= "1111111111";
                when x"C37" => data <= "1111111111";
                when x"C38" => data <= "1111111111";
                when x"C39" => data <= "1111111111";
                when x"C3A" => data <= "1111111111";
                when x"C3B" => data <= "1111111111";
                when x"C3C" => data <= "1111111111";
                when x"C3D" => data <= "1111111111";
                when x"C3E" => data <= "1111111111";
                when x"C3F" => data <= "1111111111";
                when x"C40" => data <= "1111111111";
                when x"C41" => data <= "1111111111";
                when x"C42" => data <= "1111111111";
                when x"C43" => data <= "1111111111";
                when x"C44" => data <= "1111111111";
                when x"C45" => data <= "1111111111";
                when x"C46" => data <= "1111111111";
                when x"C47" => data <= "1111111111";
                when x"C48" => data <= "1111111111";
                when x"C49" => data <= "1111111111";
                when x"C4A" => data <= "1111111111";
                when x"C4B" => data <= "1111111111";
                when x"C4C" => data <= "1111111111";
                when x"C4D" => data <= "1111111111";
                when x"C4E" => data <= "1111111111";
                when x"C4F" => data <= "1111111111";
                when x"C50" => data <= "1111111111";
                when x"C51" => data <= "1111111111";
                when x"C52" => data <= "1111111111";
                when x"C53" => data <= "1111111111";
                when x"C54" => data <= "1111111111";
                when x"C55" => data <= "1111111111";
                when x"C56" => data <= "1111111111";
                when x"C57" => data <= "1111111111";
                when x"C58" => data <= "1111111111";
                when x"C59" => data <= "1111111111";
                when x"C5A" => data <= "1111111111";
                when x"C5B" => data <= "1111111111";
                when x"C5C" => data <= "1111111111";
                when x"C5D" => data <= "1111111111";
                when x"C5E" => data <= "1111111111";
                when x"C5F" => data <= "1111111111";
                when x"C60" => data <= "1111111111";
                when x"C61" => data <= "1111111111";
                when x"C62" => data <= "1111111111";
                when x"C63" => data <= "1111111111";
                when x"C64" => data <= "1111111111";
                when x"C65" => data <= "1111111111";
                when x"C66" => data <= "1111111111";
                when x"C67" => data <= "1111111111";
                when x"C68" => data <= "1111111111";
                when x"C69" => data <= "1111111111";
                when x"C6A" => data <= "1111111111";
                when x"C6B" => data <= "1111111111";
                when x"C6C" => data <= "1111111111";
                when x"C6D" => data <= "1111111111";
                when x"C6E" => data <= "1111111111";
                when x"C6F" => data <= "1111111111";
                when x"C70" => data <= "1111111111";
                when x"C71" => data <= "1111111111";
                when x"C72" => data <= "1111111111";
                when x"C73" => data <= "1111111111";
                when x"C74" => data <= "1111111111";
                when x"C75" => data <= "1111111111";
                when x"C76" => data <= "1111111111";
                when x"C77" => data <= "1111111111";
                when x"C78" => data <= "1111111111";
                when x"C79" => data <= "1111111111";
                when x"C7A" => data <= "1111111111";
                when x"C7B" => data <= "1111111111";
                when x"C7C" => data <= "1111111111";
                when x"C7D" => data <= "1111111111";
                when x"C7E" => data <= "1111111111";
                when x"C7F" => data <= "1111111111";
                when x"C80" => data <= "1111111111";
                when x"C81" => data <= "1111111111";
                when x"C82" => data <= "1111111111";
                when x"C83" => data <= "1111111111";
                when x"C84" => data <= "1111111111";
                when x"C85" => data <= "1111111111";
                when x"C86" => data <= "1111111111";
                when x"C87" => data <= "1111111111";
                when x"C88" => data <= "1111111111";
                when x"C89" => data <= "0001111011";
                when x"C8A" => data <= "1111111111";
                when x"C8B" => data <= "1111111111";
                when x"C8C" => data <= "1111111111";
                when x"C8D" => data <= "1111111111";
                when x"C8E" => data <= "1111111111";
                when x"C8F" => data <= "1111111111";
                when x"C90" => data <= "1111111111";
                when x"C91" => data <= "1111111111";
                when x"C92" => data <= "1111111111";
                when x"C93" => data <= "1111111111";
                when x"C94" => data <= "1111111111";
                when x"C95" => data <= "1111111111";
                when x"C96" => data <= "1111111111";
                when x"C97" => data <= "1111111111";
                when x"C98" => data <= "1111111111";
                when x"C99" => data <= "1111111111";
                when x"C9A" => data <= "1111111111";
                when x"C9B" => data <= "1111111111";
                when x"C9C" => data <= "1111111111";
                when x"C9D" => data <= "1111111111";
                when x"C9E" => data <= "1111111111";
                when x"C9F" => data <= "1111111111";
                when x"CA0" => data <= "1111111111";
                when x"CA1" => data <= "1000001000";
                when x"CA2" => data <= "1111111111";
                when x"CA3" => data <= "1111111111";
                when x"CA4" => data <= "1111111111";
                when x"CA5" => data <= "1111111111";
                when x"CA6" => data <= "1111111111";
                when x"CA7" => data <= "1111111111";
                when x"CA8" => data <= "1111111111";
                when x"CA9" => data <= "1111111111";
                when x"CAA" => data <= "1111111111";
                when x"CAB" => data <= "1111111111";
                when x"CAC" => data <= "1111111111";
                when x"CAD" => data <= "1111111111";
                when x"CAE" => data <= "1111111111";
                when x"CAF" => data <= "1111111111";
                when x"CB0" => data <= "1111111111";
                when x"CB1" => data <= "1111111111";
                when x"CB2" => data <= "1111111111";
                when x"CB3" => data <= "1111111111";
                when x"CB4" => data <= "1111111111";
                when x"CB5" => data <= "1111111111";
                when x"CB6" => data <= "1111111111";
                when x"CB7" => data <= "1111111111";
                when x"CB8" => data <= "1111111111";
                when x"CB9" => data <= "1111111111";
                when x"CBA" => data <= "1111111111";
                when x"CBB" => data <= "1111111111";
                when x"CBC" => data <= "1111111111";
                when x"CBD" => data <= "1111111111";
                when x"CBE" => data <= "1111111111";
                when x"CBF" => data <= "1111111111";
                when x"CC0" => data <= "1111111111";
                when x"CC1" => data <= "1111111111";
                when x"CC2" => data <= "1111111111";
                when x"CC3" => data <= "1111111111";
                when x"CC4" => data <= "1111111111";
                when x"CC5" => data <= "1111111111";
                when x"CC6" => data <= "1111111111";
                when x"CC7" => data <= "1111111111";
                when x"CC8" => data <= "1111111111";
                when x"CC9" => data <= "1111111111";
                when x"CCA" => data <= "1111111111";
                when x"CCB" => data <= "1111111111";
                when x"CCC" => data <= "1111111111";
                when x"CCD" => data <= "1111111111";
                when x"CCE" => data <= "1111111111";
                when x"CCF" => data <= "1111111111";
                when x"CD0" => data <= "1111111111";
                when x"CD1" => data <= "1111111111";
                when x"CD2" => data <= "1111111111";
                when x"CD3" => data <= "1111111111";
                when x"CD4" => data <= "1111111111";
                when x"CD5" => data <= "1111111111";
                when x"CD6" => data <= "1111111111";
                when x"CD7" => data <= "1111111111";
                when x"CD8" => data <= "1111111111";
                when x"CD9" => data <= "1111111111";
                when x"CDA" => data <= "1111111111";
                when x"CDB" => data <= "1111111111";
                when x"CDC" => data <= "1111111111";
                when x"CDD" => data <= "1111111111";
                when x"CDE" => data <= "1111111111";
                when x"CDF" => data <= "1111111111";
                when x"CE0" => data <= "1111111111";
                when x"CE1" => data <= "1111111111";
                when x"CE2" => data <= "1111111111";
                when x"CE3" => data <= "1111111111";
                when x"CE4" => data <= "1111111111";
                when x"CE5" => data <= "1111111111";
                when x"CE6" => data <= "1111111111";
                when x"CE7" => data <= "1111111111";
                when x"CE8" => data <= "1111111111";
                when x"CE9" => data <= "1111111111";
                when x"CEA" => data <= "1111111111";
                when x"CEB" => data <= "1111111111";
                when x"CEC" => data <= "1111111111";
                when x"CED" => data <= "1111111111";
                when x"CEE" => data <= "1111111111";
                when x"CEF" => data <= "1111111111";
                when x"CF0" => data <= "1111111111";
                when x"CF1" => data <= "1111111111";
                when x"CF2" => data <= "1111111111";
                when x"CF3" => data <= "1111111111";
                when x"CF4" => data <= "1111111111";
                when x"CF5" => data <= "1111111111";
                when x"CF6" => data <= "1111111111";
                when x"CF7" => data <= "1111111111";
                when x"CF8" => data <= "1111111111";
                when x"CF9" => data <= "1111111111";
                when x"CFA" => data <= "1111111111";
                when x"CFB" => data <= "1111111111";
                when x"CFC" => data <= "1111111111";
                when x"CFD" => data <= "1111111111";
                when x"CFE" => data <= "1111111111";
                when x"CFF" => data <= "1111111111";
                when x"D00" => data <= "1111111111";
                when x"D01" => data <= "1111111111";
                when x"D02" => data <= "1111111111";
                when x"D03" => data <= "1111111111";
                when x"D04" => data <= "1111111111";
                when x"D05" => data <= "1111111111";
                when x"D06" => data <= "1111111111";
                when x"D07" => data <= "1111111111";
                when x"D08" => data <= "1111111111";
                when x"D09" => data <= "1111111111";
                when x"D0A" => data <= "1111111111";
                when x"D0B" => data <= "1111111111";
                when x"D0C" => data <= "1111111111";
                when x"D0D" => data <= "1111111111";
                when x"D0E" => data <= "1111111111";
                when x"D0F" => data <= "1111111111";
                when x"D10" => data <= "1111111111";
                when x"D11" => data <= "1111111111";
                when x"D12" => data <= "1111111111";
                when x"D13" => data <= "1111111111";
                when x"D14" => data <= "1111111111";
                when x"D15" => data <= "1111111111";
                when x"D16" => data <= "1111111111";
                when x"D17" => data <= "1111111111";
                when x"D18" => data <= "1111111111";
                when x"D19" => data <= "1111111111";
                when x"D1A" => data <= "1111111111";
                when x"D1B" => data <= "1111111111";
                when x"D1C" => data <= "1111111111";
                when x"D1D" => data <= "1111111111";
                when x"D1E" => data <= "1111111111";
                when x"D1F" => data <= "1111111111";
                when x"D20" => data <= "1111111111";
                when x"D21" => data <= "1111111111";
                when x"D22" => data <= "1111111111";
                when x"D23" => data <= "1111111111";
                when x"D24" => data <= "1111111111";
                when x"D25" => data <= "1111111111";
                when x"D26" => data <= "1111111111";
                when x"D27" => data <= "1111111111";
                when x"D28" => data <= "1111111111";
                when x"D29" => data <= "1111111111";
                when x"D2A" => data <= "1111111111";
                when x"D2B" => data <= "1111111111";
                when x"D2C" => data <= "1111111111";
                when x"D2D" => data <= "1111111111";
                when x"D2E" => data <= "1111111111";
                when x"D2F" => data <= "1111111111";
                when x"D30" => data <= "1111111111";
                when x"D31" => data <= "1111111111";
                when x"D32" => data <= "0101011000";
                when x"D33" => data <= "1111111111";
                when x"D34" => data <= "1111111111";
                when x"D35" => data <= "1111111111";
                when x"D36" => data <= "1111111111";
                when x"D37" => data <= "1111111111";
                when x"D38" => data <= "1111111111";
                when x"D39" => data <= "1111111111";
                when x"D3A" => data <= "1111111111";
                when x"D3B" => data <= "1111111111";
                when x"D3C" => data <= "1111111111";
                when x"D3D" => data <= "1111111111";
                when x"D3E" => data <= "1111111111";
                when x"D3F" => data <= "1111111111";
                when x"D40" => data <= "1111111111";
                when x"D41" => data <= "1111111111";
                when x"D42" => data <= "1111111111";
                when x"D43" => data <= "1111111111";
                when x"D44" => data <= "1111111111";
                when x"D45" => data <= "1111111111";
                when x"D46" => data <= "1111111111";
                when x"D47" => data <= "1111111111";
                when x"D48" => data <= "1111111111";
                when x"D49" => data <= "1111111111";
                when x"D4A" => data <= "1111111111";
                when x"D4B" => data <= "1111111111";
                when x"D4C" => data <= "1111111111";
                when x"D4D" => data <= "1111111111";
                when x"D4E" => data <= "1111111111";
                when x"D4F" => data <= "1111111111";
                when x"D50" => data <= "1111111111";
                when x"D51" => data <= "1111111111";
                when x"D52" => data <= "1111111111";
                when x"D53" => data <= "1111111111";
                when x"D54" => data <= "1111111111";
                when x"D55" => data <= "1111111111";
                when x"D56" => data <= "1111111111";
                when x"D57" => data <= "1111111111";
                when x"D58" => data <= "1111111111";
                when x"D59" => data <= "1111111111";
                when x"D5A" => data <= "1111111111";
                when x"D5B" => data <= "1111111111";
                when x"D5C" => data <= "1111111111";
                when x"D5D" => data <= "1111111111";
                when x"D5E" => data <= "1111111111";
                when x"D5F" => data <= "1111111111";
                when x"D60" => data <= "1111111111";
                when x"D61" => data <= "1111111111";
                when x"D62" => data <= "1111111111";
                when x"D63" => data <= "1111111111";
                when x"D64" => data <= "1111111111";
                when x"D65" => data <= "1111111111";
                when x"D66" => data <= "1111111111";
                when x"D67" => data <= "1111111111";
                when x"D68" => data <= "1111111111";
                when x"D69" => data <= "1111111111";
                when x"D6A" => data <= "1111111111";
                when x"D6B" => data <= "1111111111";
                when x"D6C" => data <= "1111111111";
                when x"D6D" => data <= "1111111111";
                when x"D6E" => data <= "1111111111";
                when x"D6F" => data <= "1111111111";
                when x"D70" => data <= "1111111111";
                when x"D71" => data <= "1111111111";
                when x"D72" => data <= "1111111111";
                when x"D73" => data <= "1111111111";
                when x"D74" => data <= "1111111111";
                when x"D75" => data <= "1111111111";
                when x"D76" => data <= "1111111111";
                when x"D77" => data <= "1111111111";
                when x"D78" => data <= "1111111111";
                when x"D79" => data <= "1111111111";
                when x"D7A" => data <= "1111111111";
                when x"D7B" => data <= "1111111111";
                when x"D7C" => data <= "1111111111";
                when x"D7D" => data <= "1111111111";
                when x"D7E" => data <= "1111111111";
                when x"D7F" => data <= "1111111111";
                when x"D80" => data <= "1111111111";
                when x"D81" => data <= "1111111111";
                when x"D82" => data <= "1111111111";
                when x"D83" => data <= "1111111111";
                when x"D84" => data <= "1111111111";
                when x"D85" => data <= "1111111111";
                when x"D86" => data <= "1111111111";
                when x"D87" => data <= "1111111111";
                when x"D88" => data <= "1111111111";
                when x"D89" => data <= "1111111111";
                when x"D8A" => data <= "1111111111";
                when x"D8B" => data <= "1111111111";
                when x"D8C" => data <= "1111111111";
                when x"D8D" => data <= "1111111111";
                when x"D8E" => data <= "1111111111";
                when x"D8F" => data <= "1111111111";
                when x"D90" => data <= "1111111111";
                when x"D91" => data <= "1111111111";
                when x"D92" => data <= "1111111111";
                when x"D93" => data <= "1111111111";
                when x"D94" => data <= "1111111111";
                when x"D95" => data <= "1111111111";
                when x"D96" => data <= "1111111111";
                when x"D97" => data <= "1111111111";
                when x"D98" => data <= "1111111111";
                when x"D99" => data <= "1111111111";
                when x"D9A" => data <= "1111111111";
                when x"D9B" => data <= "1111111111";
                when x"D9C" => data <= "1111111111";
                when x"D9D" => data <= "1111111111";
                when x"D9E" => data <= "1111111111";
                when x"D9F" => data <= "1111111111";
                when x"DA0" => data <= "1111111111";
                when x"DA1" => data <= "1111111111";
                when x"DA2" => data <= "1111111111";
                when x"DA3" => data <= "1111111111";
                when x"DA4" => data <= "1111111111";
                when x"DA5" => data <= "1111111111";
                when x"DA6" => data <= "1111111111";
                when x"DA7" => data <= "1111111111";
                when x"DA8" => data <= "1111111111";
                when x"DA9" => data <= "1111111111";
                when x"DAA" => data <= "1111111111";
                when x"DAB" => data <= "1111111111";
                when x"DAC" => data <= "1111111111";
                when x"DAD" => data <= "1111111111";
                when x"DAE" => data <= "1111111111";
                when x"DAF" => data <= "1111111111";
                when x"DB0" => data <= "1111111111";
                when x"DB1" => data <= "1111111111";
                when x"DB2" => data <= "1111111111";
                when x"DB3" => data <= "1111111111";
                when x"DB4" => data <= "1111111111";
                when x"DB5" => data <= "1111111111";
                when x"DB6" => data <= "1111111111";
                when x"DB7" => data <= "1111111111";
                when x"DB8" => data <= "1111111111";
                when x"DB9" => data <= "1111111111";
                when x"DBA" => data <= "1111111111";
                when x"DBB" => data <= "1111111111";
                when x"DBC" => data <= "1111111111";
                when x"DBD" => data <= "1111111111";
                when x"DBE" => data <= "1111111111";
                when x"DBF" => data <= "1111111111";
                when x"DC0" => data <= "1111111111";
                when x"DC1" => data <= "1111111111";
                when x"DC2" => data <= "1111111111";
                when x"DC3" => data <= "1111111111";
                when x"DC4" => data <= "1111111111";
                when x"DC5" => data <= "1111111111";
                when x"DC6" => data <= "1111111111";
                when x"DC7" => data <= "1111111111";
                when x"DC8" => data <= "1111111111";
                when x"DC9" => data <= "1111111111";
                when x"DCA" => data <= "1111111111";
                when x"DCB" => data <= "1111111111";
                when x"DCC" => data <= "1111111111";
                when x"DCD" => data <= "1111111111";
                when x"DCE" => data <= "1111111111";
                when x"DCF" => data <= "1111111111";
                when x"DD0" => data <= "1111111111";
                when x"DD1" => data <= "1111111111";
                when x"DD2" => data <= "1000001000";
                when x"DD3" => data <= "1111111111";
                when x"DD4" => data <= "1111111111";
                when x"DD5" => data <= "1111111111";
                when x"DD6" => data <= "1111111111";
                when x"DD7" => data <= "1111111111";
                when x"DD8" => data <= "1111111111";
                when x"DD9" => data <= "1111111111";
                when x"DDA" => data <= "1111111111";
                when x"DDB" => data <= "1111111111";
                when x"DDC" => data <= "1111111111";
                when x"DDD" => data <= "1111111111";
                when x"DDE" => data <= "1111111111";
                when x"DDF" => data <= "1111111111";
                when x"DE0" => data <= "1111111111";
                when x"DE1" => data <= "1111111111";
                when x"DE2" => data <= "1111111111";
                when x"DE3" => data <= "1000111101";
                when x"DE4" => data <= "1111111111";
                when x"DE5" => data <= "1111111111";
                when x"DE6" => data <= "1111111111";
                when x"DE7" => data <= "1111111111";
                when x"DE8" => data <= "1111111111";
                when x"DE9" => data <= "1111111111";
                when x"DEA" => data <= "1111111111";
                when x"DEB" => data <= "1111111111";
                when x"DEC" => data <= "1111111111";
                when x"DED" => data <= "1111111111";
                when x"DEE" => data <= "1111111111";
                when x"DEF" => data <= "1111111111";
                when x"DF0" => data <= "1111111111";
                when x"DF1" => data <= "1111111111";
                when x"DF2" => data <= "1111111111";
                when x"DF3" => data <= "1111111111";
                when x"DF4" => data <= "1111111111";
                when x"DF5" => data <= "1111111111";
                when x"DF6" => data <= "1111111111";
                when x"DF7" => data <= "1111111111";
                when x"DF8" => data <= "1111111111";
                when x"DF9" => data <= "1111111111";
                when x"DFA" => data <= "1111111111";
                when x"DFB" => data <= "1111111111";
                when x"DFC" => data <= "1111111111";
                when x"DFD" => data <= "1111111111";
                when x"DFE" => data <= "1111111111";
                when x"DFF" => data <= "1111111111";
                when x"E00" => data <= "1111111111";
                when x"E01" => data <= "1111111111";
                when x"E02" => data <= "1111111111";
                when x"E03" => data <= "1111111111";
                when x"E04" => data <= "1111111111";
                when x"E05" => data <= "1111111111";
                when x"E06" => data <= "1111111111";
                when x"E07" => data <= "1111111111";
                when x"E08" => data <= "1111111111";
                when x"E09" => data <= "1111111111";
                when x"E0A" => data <= "1111111111";
                when x"E0B" => data <= "1111111111";
                when x"E0C" => data <= "1111111111";
                when x"E0D" => data <= "1111111111";
                when x"E0E" => data <= "1111111111";
                when x"E0F" => data <= "1111111111";
                when x"E10" => data <= "1111111111";
                when x"E11" => data <= "1111111111";
                when x"E12" => data <= "1111111111";
                when x"E13" => data <= "1111111111";
                when x"E14" => data <= "1111111111";
                when x"E15" => data <= "1111111111";
                when x"E16" => data <= "1111111111";
                when x"E17" => data <= "1111111111";
                when x"E18" => data <= "1111111111";
                when x"E19" => data <= "1111111111";
                when x"E1A" => data <= "1111111111";
                when x"E1B" => data <= "1111111111";
                when x"E1C" => data <= "1111111111";
                when x"E1D" => data <= "1111111111";
                when x"E1E" => data <= "1111111111";
                when x"E1F" => data <= "1111111111";
                when x"E20" => data <= "1111111111";
                when x"E21" => data <= "0000100100";
                when x"E22" => data <= "1111111111";
                when x"E23" => data <= "1111111111";
                when x"E24" => data <= "1111111111";
                when x"E25" => data <= "1111111111";
                when x"E26" => data <= "1111111111";
                when x"E27" => data <= "1111111111";
                when x"E28" => data <= "1111111111";
                when x"E29" => data <= "1111111111";
                when x"E2A" => data <= "1111111111";
                when x"E2B" => data <= "1111111111";
                when x"E2C" => data <= "1111111111";
                when x"E2D" => data <= "1111111111";
                when x"E2E" => data <= "1111111111";
                when x"E2F" => data <= "1111111111";
                when x"E30" => data <= "1111111111";
                when x"E31" => data <= "1111111111";
                when x"E32" => data <= "1111111111";
                when x"E33" => data <= "1111111111";
                when x"E34" => data <= "1111111111";
                when x"E35" => data <= "1000001000";
                when x"E36" => data <= "1111111111";
                when x"E37" => data <= "1111111111";
                when x"E38" => data <= "1111111111";
                when x"E39" => data <= "1111111111";
                when x"E3A" => data <= "1111111111";
                when x"E3B" => data <= "1111111111";
                when x"E3C" => data <= "1111111111";
                when x"E3D" => data <= "1111111111";
                when x"E3E" => data <= "1111111111";
                when x"E3F" => data <= "1111111111";
                when x"E40" => data <= "1111111111";
                when x"E41" => data <= "1111111111";
                when x"E42" => data <= "1111111111";
                when x"E43" => data <= "1111111111";
                when x"E44" => data <= "1111111111";
                when x"E45" => data <= "1111111111";
                when x"E46" => data <= "1111111111";
                when x"E47" => data <= "1111111111";
                when x"E48" => data <= "1111111111";
                when x"E49" => data <= "1111111111";
                when x"E4A" => data <= "1111111111";
                when x"E4B" => data <= "1111111111";
                when x"E4C" => data <= "1111111111";
                when x"E4D" => data <= "1111111111";
                when x"E4E" => data <= "1111111111";
                when x"E4F" => data <= "1111111111";
                when x"E50" => data <= "1111111111";
                when x"E51" => data <= "1111111111";
                when x"E52" => data <= "1111111111";
                when x"E53" => data <= "1111111111";
                when x"E54" => data <= "1111111111";
                when x"E55" => data <= "1111111111";
                when x"E56" => data <= "1111111111";
                when x"E57" => data <= "1111111111";
                when x"E58" => data <= "1111111111";
                when x"E59" => data <= "1111111111";
                when x"E5A" => data <= "1111111111";
                when x"E5B" => data <= "1111111111";
                when x"E5C" => data <= "1111111111";
                when x"E5D" => data <= "1111111111";
                when x"E5E" => data <= "1111111111";
                when x"E5F" => data <= "1111111111";
                when x"E60" => data <= "1111111111";
                when x"E61" => data <= "1111111111";
                when x"E62" => data <= "1111111111";
                when x"E63" => data <= "1111111111";
                when x"E64" => data <= "1111111111";
                when x"E65" => data <= "1111111111";
                when x"E66" => data <= "1111111111";
                when x"E67" => data <= "1111111111";
                when x"E68" => data <= "1111111111";
                when x"E69" => data <= "1111111111";
                when x"E6A" => data <= "1111111111";
                when x"E6B" => data <= "1111111111";
                when x"E6C" => data <= "1111111111";
                when x"E6D" => data <= "1111111111";
                when x"E6E" => data <= "1111111111";
                when x"E6F" => data <= "1111111111";
                when x"E70" => data <= "1111111111";
                when x"E71" => data <= "1111111111";
                when x"E72" => data <= "1111111111";
                when x"E73" => data <= "1111111111";
                when x"E74" => data <= "1111111111";
                when x"E75" => data <= "1111111111";
                when x"E76" => data <= "1111111111";
                when x"E77" => data <= "1111111111";
                when x"E78" => data <= "1111111111";
                when x"E79" => data <= "1111111111";
                when x"E7A" => data <= "1111111111";
                when x"E7B" => data <= "0110001100";
                when x"E7C" => data <= "1111111111";
                when x"E7D" => data <= "1111111111";
                when x"E7E" => data <= "1111111111";
                when x"E7F" => data <= "1111111111";
                when x"E80" => data <= "1111111111";
                when x"E81" => data <= "1111111111";
                when x"E82" => data <= "1111111111";
                when x"E83" => data <= "1111111111";
                when x"E84" => data <= "1111111111";
                when x"E85" => data <= "1111111111";
                when x"E86" => data <= "1111111111";
                when x"E87" => data <= "1111111111";
                when x"E88" => data <= "1111111111";
                when x"E89" => data <= "1111111111";
                when x"E8A" => data <= "1111111111";
                when x"E8B" => data <= "1111111111";
                when x"E8C" => data <= "1111111111";
                when x"E8D" => data <= "1111111111";
                when x"E8E" => data <= "1111111111";
                when x"E8F" => data <= "1111111111";
                when x"E90" => data <= "1111111111";
                when x"E91" => data <= "1111111111";
                when x"E92" => data <= "1111111111";
                when x"E93" => data <= "1111111111";
                when x"E94" => data <= "1111111111";
                when x"E95" => data <= "1111111111";
                when x"E96" => data <= "1111111111";
                when x"E97" => data <= "1111111111";
                when x"E98" => data <= "1111111111";
                when x"E99" => data <= "1111111111";
                when x"E9A" => data <= "1111111111";
                when x"E9B" => data <= "1111111111";
                when x"E9C" => data <= "1111111111";
                when x"E9D" => data <= "1111111111";
                when x"E9E" => data <= "1111111111";
                when x"E9F" => data <= "1111111111";
                when x"EA0" => data <= "1111111111";
                when x"EA1" => data <= "1111111111";
                when x"EA2" => data <= "1111111111";
                when x"EA3" => data <= "1111111111";
                when x"EA4" => data <= "1111111111";
                when x"EA5" => data <= "1111111111";
                when x"EA6" => data <= "1111111111";
                when x"EA7" => data <= "1111111111";
                when x"EA8" => data <= "1111111111";
                when x"EA9" => data <= "1111111111";
                when x"EAA" => data <= "1111111111";
                when x"EAB" => data <= "1111111111";
                when x"EAC" => data <= "1111111111";
                when x"EAD" => data <= "1111111111";
                when x"EAE" => data <= "1111111111";
                when x"EAF" => data <= "1111111111";
                when x"EB0" => data <= "1111111111";
                when x"EB1" => data <= "1111111111";
                when x"EB2" => data <= "1111111111";
                when x"EB3" => data <= "1111111111";
                when x"EB4" => data <= "1111111111";
                when x"EB5" => data <= "1000001000";
                when x"EB6" => data <= "1111111111";
                when x"EB7" => data <= "1111111111";
                when x"EB8" => data <= "1111111111";
                when x"EB9" => data <= "1111111111";
                when x"EBA" => data <= "1111111111";
                when x"EBB" => data <= "1111111111";
                when x"EBC" => data <= "1111111111";
                when x"EBD" => data <= "1111111111";
                when x"EBE" => data <= "1111111111";
                when x"EBF" => data <= "1111111111";
                when x"EC0" => data <= "1111111111";
                when x"EC1" => data <= "1111111111";
                when x"EC2" => data <= "1111111111";
                when x"EC3" => data <= "1111111111";
                when x"EC4" => data <= "1111111111";
                when x"EC5" => data <= "1111111111";
                when x"EC6" => data <= "1111111111";
                when x"EC7" => data <= "1111111111";
                when x"EC8" => data <= "1111111111";
                when x"EC9" => data <= "1111111111";
                when x"ECA" => data <= "1111111111";
                when x"ECB" => data <= "1111111111";
                when x"ECC" => data <= "1111111111";
                when x"ECD" => data <= "1111111111";
                when x"ECE" => data <= "1111111111";
                when x"ECF" => data <= "1111111111";
                when x"ED0" => data <= "1111111111";
                when x"ED1" => data <= "1111111111";
                when x"ED2" => data <= "1111111111";
                when x"ED3" => data <= "1111111111";
                when x"ED4" => data <= "1111111111";
                when x"ED5" => data <= "1111111111";
                when x"ED6" => data <= "1111111111";
                when x"ED7" => data <= "1111111111";
                when x"ED8" => data <= "1111111111";
                when x"ED9" => data <= "1111111111";
                when x"EDA" => data <= "1111111111";
                when x"EDB" => data <= "1111111111";
                when x"EDC" => data <= "1111111111";
                when x"EDD" => data <= "1111111111";
                when x"EDE" => data <= "1111111111";
                when x"EDF" => data <= "1111111111";
                when x"EE0" => data <= "1111111111";
                when x"EE1" => data <= "1111111111";
                when x"EE2" => data <= "1111111111";
                when x"EE3" => data <= "1111111111";
                when x"EE4" => data <= "1111111111";
                when x"EE5" => data <= "1111111111";
                when x"EE6" => data <= "1111111111";
                when x"EE7" => data <= "1111111111";
                when x"EE8" => data <= "1111111111";
                when x"EE9" => data <= "1111111111";
                when x"EEA" => data <= "1111111111";
                when x"EEB" => data <= "1111111111";
                when x"EEC" => data <= "1111111111";
                when x"EED" => data <= "1111111111";
                when x"EEE" => data <= "1111111111";
                when x"EEF" => data <= "1111111111";
                when x"EF0" => data <= "1111111111";
                when x"EF1" => data <= "1111111111";
                when x"EF2" => data <= "1111111111";
                when x"EF3" => data <= "1111111111";
                when x"EF4" => data <= "1111111111";
                when x"EF5" => data <= "1111111111";
                when x"EF6" => data <= "1111111111";
                when x"EF7" => data <= "1111111111";
                when x"EF8" => data <= "1111111111";
                when x"EF9" => data <= "1111111111";
                when x"EFA" => data <= "1111111111";
                when x"EFB" => data <= "1111111111";
                when x"EFC" => data <= "1111111111";
                when x"EFD" => data <= "1111111111";
                when x"EFE" => data <= "1111111111";
                when x"EFF" => data <= "1111111111";
                when x"F00" => data <= "1111111111";
                when x"F01" => data <= "1111111111";
                when x"F02" => data <= "1111111111";
                when x"F03" => data <= "1111111111";
                when x"F04" => data <= "1111111111";
                when x"F05" => data <= "1111111111";
                when x"F06" => data <= "1111111111";
                when x"F07" => data <= "1111111111";
                when x"F08" => data <= "1111111111";
                when x"F09" => data <= "1000001000";
                when x"F0A" => data <= "1111111111";
                when x"F0B" => data <= "1111111111";
                when x"F0C" => data <= "1111111111";
                when x"F0D" => data <= "1111111111";
                when x"F0E" => data <= "1111111111";
                when x"F0F" => data <= "1111111111";
                when x"F10" => data <= "1111111111";
                when x"F11" => data <= "1111111111";
                when x"F12" => data <= "1111111111";
                when x"F13" => data <= "1111111111";
                when x"F14" => data <= "1111111111";
                when x"F15" => data <= "1111111111";
                when x"F16" => data <= "1111111111";
                when x"F17" => data <= "1111111111";
                when x"F18" => data <= "1111111111";
                when x"F19" => data <= "1111111111";
                when x"F1A" => data <= "1111111111";
                when x"F1B" => data <= "1111111111";
                when x"F1C" => data <= "1111111111";
                when x"F1D" => data <= "1111111111";
                when x"F1E" => data <= "1111111111";
                when x"F1F" => data <= "1111111111";
                when x"F20" => data <= "1111111111";
                when x"F21" => data <= "1111111111";
                when x"F22" => data <= "1111111111";
                when x"F23" => data <= "1111111111";
                when x"F24" => data <= "1111111111";
                when x"F25" => data <= "1111111111";
                when x"F26" => data <= "1111111111";
                when x"F27" => data <= "1111111111";
                when x"F28" => data <= "1111111111";
                when x"F29" => data <= "1111111111";
                when x"F2A" => data <= "1111111111";
                when x"F2B" => data <= "1111111111";
                when x"F2C" => data <= "1111111111";
                when x"F2D" => data <= "1111111111";
                when x"F2E" => data <= "1111111111";
                when x"F2F" => data <= "1111111111";
                when x"F30" => data <= "1111111111";
                when x"F31" => data <= "1111111111";
                when x"F32" => data <= "1111111111";
                when x"F33" => data <= "1111111111";
                when x"F34" => data <= "1000001000";
                when x"F35" => data <= "1111111111";
                when x"F36" => data <= "1111111111";
                when x"F37" => data <= "1111111111";
                when x"F38" => data <= "1111111111";
                when x"F39" => data <= "1111111111";
                when x"F3A" => data <= "1111111111";
                when x"F3B" => data <= "1111111111";
                when x"F3C" => data <= "1111111111";
                when x"F3D" => data <= "1111111111";
                when x"F3E" => data <= "1111111111";
                when x"F3F" => data <= "1111111111";
                when x"F40" => data <= "1111111111";
                when x"F41" => data <= "1111111111";
                when x"F42" => data <= "1111111111";
                when x"F43" => data <= "1111111111";
                when x"F44" => data <= "1111111111";
                when x"F45" => data <= "1111111111";
                when x"F46" => data <= "1111111111";
                when x"F47" => data <= "1111111111";
                when x"F48" => data <= "1111111111";
                when x"F49" => data <= "1111111111";
                when x"F4A" => data <= "1111111111";
                when x"F4B" => data <= "1111111111";
                when x"F4C" => data <= "1111111111";
                when x"F4D" => data <= "1111111111";
                when x"F4E" => data <= "1111111111";
                when x"F4F" => data <= "1111111111";
                when x"F50" => data <= "1111111111";
                when x"F51" => data <= "1111111111";
                when x"F52" => data <= "1111111111";
                when x"F53" => data <= "1111111111";
                when x"F54" => data <= "1111111111";
                when x"F55" => data <= "1111111111";
                when x"F56" => data <= "1111111111";
                when x"F57" => data <= "1111111111";
                when x"F58" => data <= "1111111111";
                when x"F59" => data <= "1111111111";
                when x"F5A" => data <= "1111111111";
                when x"F5B" => data <= "1111111111";
                when x"F5C" => data <= "1111111111";
                when x"F5D" => data <= "1111111111";
                when x"F5E" => data <= "1111111111";
                when x"F5F" => data <= "1111111111";
                when x"F60" => data <= "1111111111";
                when x"F61" => data <= "1111111111";
                when x"F62" => data <= "1000001000";
                when x"F63" => data <= "1111111111";
                when x"F64" => data <= "1111111111";
                when x"F65" => data <= "1111111111";
                when x"F66" => data <= "1111111111";
                when x"F67" => data <= "1111111111";
                when x"F68" => data <= "1111111111";
                when x"F69" => data <= "1111111111";
                when x"F6A" => data <= "1111111111";
                when x"F6B" => data <= "1111111111";
                when x"F6C" => data <= "1111111111";
                when x"F6D" => data <= "1111111111";
                when x"F6E" => data <= "1111111111";
                when x"F6F" => data <= "1111111111";
                when x"F70" => data <= "1111111111";
                when x"F71" => data <= "1111111111";
                when x"F72" => data <= "1111111111";
                when x"F73" => data <= "1111111111";
                when x"F74" => data <= "1111111111";
                when x"F75" => data <= "1111111111";
                when x"F76" => data <= "1111111111";
                when x"F77" => data <= "1111111111";
                when x"F78" => data <= "1111111111";
                when x"F79" => data <= "1111111111";
                when x"F7A" => data <= "1111111111";
                when x"F7B" => data <= "1111111111";
                when x"F7C" => data <= "1111111111";
                when x"F7D" => data <= "1111111111";
                when x"F7E" => data <= "1111111111";
                when x"F7F" => data <= "1111111111";
                when x"F80" => data <= "1111111111";
                when x"F81" => data <= "1111111111";
                when x"F82" => data <= "1111111111";
                when x"F83" => data <= "1111111111";
                when x"F84" => data <= "1111111111";
                when x"F85" => data <= "1111111111";
                when x"F86" => data <= "1111111111";
                when x"F87" => data <= "1111111111";
                when x"F88" => data <= "1111111111";
                when x"F89" => data <= "1111111111";
                when x"F8A" => data <= "1111111111";
                when x"F8B" => data <= "1111111111";
                when x"F8C" => data <= "1111111111";
                when x"F8D" => data <= "1111111111";
                when x"F8E" => data <= "1111111111";
                when x"F8F" => data <= "1111111111";
                when x"F90" => data <= "1111111111";
                when x"F91" => data <= "1111111111";
                when x"F92" => data <= "1111111111";
                when x"F93" => data <= "1111111111";
                when x"F94" => data <= "1111111111";
                when x"F95" => data <= "1111111111";
                when x"F96" => data <= "1111111111";
                when x"F97" => data <= "1111111111";
                when x"F98" => data <= "1111111111";
                when x"F99" => data <= "1111111111";
                when x"F9A" => data <= "1111111111";
                when x"F9B" => data <= "1111111111";
                when x"F9C" => data <= "1111111111";
                when x"F9D" => data <= "1111111111";
                when x"F9E" => data <= "1111111111";
                when x"F9F" => data <= "1111111111";
                when x"FA0" => data <= "1111111111";
                when x"FA1" => data <= "1111111111";
                when x"FA2" => data <= "1111111111";
                when x"FA3" => data <= "1111111111";
                when x"FA4" => data <= "1111111111";
                when x"FA5" => data <= "1111111111";
                when x"FA6" => data <= "1111111111";
                when x"FA7" => data <= "1111111111";
                when x"FA8" => data <= "1111111111";
                when x"FA9" => data <= "1111111111";
                when x"FAA" => data <= "1111111111";
                when x"FAB" => data <= "1111111111";
                when x"FAC" => data <= "1111111111";
                when x"FAD" => data <= "1111111111";
                when x"FAE" => data <= "1111111111";
                when x"FAF" => data <= "1111111111";
                when x"FB0" => data <= "1111111111";
                when x"FB1" => data <= "1111111111";
                when x"FB2" => data <= "1111111111";
                when x"FB3" => data <= "1111111111";
                when x"FB4" => data <= "1111111111";
                when x"FB5" => data <= "1111111111";
                when x"FB6" => data <= "1111111111";
                when x"FB7" => data <= "1111111111";
                when x"FB8" => data <= "1111111111";
                when x"FB9" => data <= "1111111111";
                when x"FBA" => data <= "0100000111";
                when x"FBB" => data <= "1111111111";
                when x"FBC" => data <= "1111111111";
                when x"FBD" => data <= "1111111111";
                when x"FBE" => data <= "1000001000";
                when x"FBF" => data <= "1111111111";
                when x"FC0" => data <= "1111111111";
                when x"FC1" => data <= "1111111111";
                when x"FC2" => data <= "1111111111";
                when x"FC3" => data <= "1111111111";
                when x"FC4" => data <= "1111111111";
                when x"FC5" => data <= "1111111111";
                when x"FC6" => data <= "1111111111";
                when x"FC7" => data <= "1111111111";
                when x"FC8" => data <= "1111111111";
                when x"FC9" => data <= "1111111111";
                when x"FCA" => data <= "1111111111";
                when x"FCB" => data <= "1111111111";
                when x"FCC" => data <= "1111111111";
                when x"FCD" => data <= "1111111111";
                when x"FCE" => data <= "1111111111";
                when x"FCF" => data <= "1111111111";
                when x"FD0" => data <= "1111111111";
                when x"FD1" => data <= "1111111111";
                when x"FD2" => data <= "1111111111";
                when x"FD3" => data <= "1111111111";
                when x"FD4" => data <= "1111111111";
                when x"FD5" => data <= "1111111111";
                when x"FD6" => data <= "1111111111";
                when x"FD7" => data <= "1111111111";
                when x"FD8" => data <= "1111111111";
                when x"FD9" => data <= "1111111111";
                when x"FDA" => data <= "1111111111";
                when x"FDB" => data <= "1111111111";
                when x"FDC" => data <= "1111111111";
                when x"FDD" => data <= "1111111111";
                when x"FDE" => data <= "1111111111";
                when x"FDF" => data <= "1111111111";
                when x"FE0" => data <= "1111111111";
                when x"FE1" => data <= "1111111111";
                when x"FE2" => data <= "1111111111";
                when x"FE3" => data <= "1111111111";
                when x"FE4" => data <= "1111111111";
                when x"FE5" => data <= "1111111111";
                when x"FE6" => data <= "1111111111";
                when x"FE7" => data <= "1111111111";
                when x"FE8" => data <= "1111111111";
                when x"FE9" => data <= "1111111111";
                when x"FEA" => data <= "1111111111";
                when x"FEB" => data <= "1111111111";
                when x"FEC" => data <= "1111111111";
                when x"FED" => data <= "1111111111";
                when x"FEE" => data <= "1111111111";
                when x"FEF" => data <= "1111111111";
                when x"FF0" => data <= "1111111111";
                when x"FF1" => data <= "1111111111";
                when x"FF2" => data <= "1111111111";
                when x"FF3" => data <= "1111111111";
                when x"FF4" => data <= "1111111111";
                when x"FF5" => data <= "1111111111";
                when x"FF6" => data <= "1111111111";
                when x"FF7" => data <= "1111111111";
                when x"FF8" => data <= "1111111111";
                when x"FF9" => data <= "1111111111";
                when x"FFA" => data <= "1111111111";
                when x"FFB" => data <= "1111111111";
                when x"FFC" => data <= "1111111111";
                when x"FFD" => data <= "1111111111";
                when x"FFE" => data <= "1111111111";
                when x"FFF" => data <= "1111111111";
                when x"1000" => data <= "1111111111";
                when x"1001" => data <= "1111111111";
                when x"1002" => data <= "1111111111";
                when x"1003" => data <= "1111111111";
                when x"1004" => data <= "1111111111";
                when x"1005" => data <= "1111111111";
                when x"1006" => data <= "1111111111";
                when x"1007" => data <= "1111111111";
                when x"1008" => data <= "1111111111";
                when x"1009" => data <= "1111111111";
                when x"100A" => data <= "1111111111";
                when x"100B" => data <= "1111111111";
                when x"100C" => data <= "1111111111";
                when x"100D" => data <= "1111111111";
                when x"100E" => data <= "1111111111";
                when x"100F" => data <= "1111111111";
                when x"1010" => data <= "1111111111";
                when x"1011" => data <= "1111111111";
                when x"1012" => data <= "1111111111";
                when x"1013" => data <= "1111111111";
                when x"1014" => data <= "1111111111";
                when x"1015" => data <= "1111111111";
                when x"1016" => data <= "1111111111";
                when x"1017" => data <= "1111111111";
                when x"1018" => data <= "1111111111";
                when x"1019" => data <= "1111111111";
                when x"101A" => data <= "1111111111";
                when x"101B" => data <= "1111111111";
                when x"101C" => data <= "1111111111";
                when x"101D" => data <= "1111111111";
                when x"101E" => data <= "1111111111";
                when x"101F" => data <= "1111111111";
                when x"1020" => data <= "1111111111";
                when x"1021" => data <= "1111111111";
                when x"1022" => data <= "1111111111";
                when x"1023" => data <= "1111111111";
                when x"1024" => data <= "1111111111";
                when x"1025" => data <= "1111111111";
                when x"1026" => data <= "1111111111";
                when x"1027" => data <= "1111111111";
                when x"1028" => data <= "1111111111";
                when x"1029" => data <= "1111111111";
                when x"102A" => data <= "1111111111";
                when x"102B" => data <= "1111111111";
                when x"102C" => data <= "1111111111";
                when x"102D" => data <= "1111111111";
                when x"102E" => data <= "1111111111";
                when x"102F" => data <= "1111111111";
                when x"1030" => data <= "1111111111";
                when x"1031" => data <= "1111111111";
                when x"1032" => data <= "1111111111";
                when x"1033" => data <= "1111111111";
                when x"1034" => data <= "1111111111";
                when x"1035" => data <= "1111111111";
                when x"1036" => data <= "1111111111";
                when x"1037" => data <= "1111111111";
                when x"1038" => data <= "1111111111";
                when x"1039" => data <= "1111111111";
                when x"103A" => data <= "1111111111";
                when x"103B" => data <= "1111111111";
                when x"103C" => data <= "1111111111";
                when x"103D" => data <= "1111111111";
                when x"103E" => data <= "1111111111";
                when x"103F" => data <= "1111111111";
                when x"1040" => data <= "1111111111";
                when x"1041" => data <= "1111111111";
                when x"1042" => data <= "1111111111";
                when x"1043" => data <= "1111111111";
                when x"1044" => data <= "1111111111";
                when x"1045" => data <= "1111111111";
                when x"1046" => data <= "1111111111";
                when x"1047" => data <= "1111111111";
                when x"1048" => data <= "1111111111";
                when x"1049" => data <= "1111111111";
                when x"104A" => data <= "1111111111";
                when x"104B" => data <= "1111111111";
                when x"104C" => data <= "1111111111";
                when x"104D" => data <= "1111111111";
                when x"104E" => data <= "1111111111";
                when x"104F" => data <= "1111111111";
                when x"1050" => data <= "1111111111";
                when x"1051" => data <= "1111111111";
                when x"1052" => data <= "1111111111";
                when x"1053" => data <= "1111111111";
                when x"1054" => data <= "1111111111";
                when x"1055" => data <= "1111111111";
                when x"1056" => data <= "1111111111";
                when x"1057" => data <= "1111111111";
                when x"1058" => data <= "1111111111";
                when x"1059" => data <= "1111111111";
                when x"105A" => data <= "1111111111";
                when x"105B" => data <= "1111111111";
                when x"105C" => data <= "1111111111";
                when x"105D" => data <= "1111111111";
                when x"105E" => data <= "1111111111";
                when x"105F" => data <= "1111111111";
                when x"1060" => data <= "1111111111";
                when x"1061" => data <= "1111111111";
                when x"1062" => data <= "1111111111";
                when x"1063" => data <= "1111111111";
                when x"1064" => data <= "1111111111";
                when x"1065" => data <= "1111111111";
                when x"1066" => data <= "1111111111";
                when x"1067" => data <= "1111111111";
                when x"1068" => data <= "1111111111";
                when x"1069" => data <= "1111111111";
                when x"106A" => data <= "1111111111";
                when x"106B" => data <= "1111111111";
                when x"106C" => data <= "1111111111";
                when x"106D" => data <= "1111111111";
                when x"106E" => data <= "1111111111";
                when x"106F" => data <= "1111111111";
                when x"1070" => data <= "1111111111";
                when x"1071" => data <= "1111111111";
                when x"1072" => data <= "1111111111";
                when x"1073" => data <= "1111111111";
                when x"1074" => data <= "1111111111";
                when x"1075" => data <= "1111111111";
                when x"1076" => data <= "1111111111";
                when x"1077" => data <= "1111111111";
                when x"1078" => data <= "1111111111";
                when x"1079" => data <= "1111111111";
                when x"107A" => data <= "1111111111";
                when x"107B" => data <= "1111111111";
                when x"107C" => data <= "1111111111";
                when x"107D" => data <= "1111111111";
                when x"107E" => data <= "1111111111";
                when x"107F" => data <= "1111111111";
                when x"1080" => data <= "1111111111";
                when x"1081" => data <= "1111111111";
                when x"1082" => data <= "1111111111";
                when x"1083" => data <= "1111111111";
                when x"1084" => data <= "1111111111";
                when x"1085" => data <= "1111111111";
                when x"1086" => data <= "1111111111";
                when x"1087" => data <= "1111111111";
                when x"1088" => data <= "1111111111";
                when x"1089" => data <= "1111111111";
                when x"108A" => data <= "1111111111";
                when x"108B" => data <= "1111111111";
                when x"108C" => data <= "1111111111";
                when x"108D" => data <= "1111111111";
                when x"108E" => data <= "1111111111";
                when x"108F" => data <= "1111111111";
                when x"1090" => data <= "1111111111";
                when x"1091" => data <= "1000001000";
                when x"1092" => data <= "1111111111";
                when x"1093" => data <= "1111111111";
                when x"1094" => data <= "1111111111";
                when x"1095" => data <= "1111111111";
                when x"1096" => data <= "1111111111";
                when x"1097" => data <= "1111111111";
                when x"1098" => data <= "1000001000";
                when x"1099" => data <= "1111111111";
                when x"109A" => data <= "1111111111";
                when x"109B" => data <= "1111111111";
                when x"109C" => data <= "1111111111";
                when x"109D" => data <= "1111111111";
                when x"109E" => data <= "1111111111";
                when x"109F" => data <= "1111111111";
                when x"10A0" => data <= "1111111111";
                when x"10A1" => data <= "1111111111";
                when x"10A2" => data <= "1111111111";
                when x"10A3" => data <= "1111111111";
                when x"10A4" => data <= "1111111111";
                when x"10A5" => data <= "1111111111";
                when x"10A6" => data <= "1111111111";
                when x"10A7" => data <= "1111111111";
                when x"10A8" => data <= "1111111111";
                when x"10A9" => data <= "1111111111";
                when x"10AA" => data <= "1111111111";
                when x"10AB" => data <= "1011011100";
                when x"10AC" => data <= "1111111111";
                when x"10AD" => data <= "1111111111";
                when x"10AE" => data <= "1111111111";
                when x"10AF" => data <= "1111111111";
                when x"10B0" => data <= "1111111111";
                when x"10B1" => data <= "1111111111";
                when x"10B2" => data <= "1111111111";
                when x"10B3" => data <= "1111111111";
                when x"10B4" => data <= "1111111111";
                when x"10B5" => data <= "1111111111";
                when x"10B6" => data <= "1111111111";
                when x"10B7" => data <= "1111111111";
                when x"10B8" => data <= "1111111111";
                when x"10B9" => data <= "1111111111";
                when x"10BA" => data <= "1111111111";
                when x"10BB" => data <= "1111111111";
                when x"10BC" => data <= "1111111111";
                when x"10BD" => data <= "1111111111";
                when x"10BE" => data <= "1111111111";
                when x"10BF" => data <= "1111111111";
                when x"10C0" => data <= "1111111111";
                when x"10C1" => data <= "1111111111";
                when x"10C2" => data <= "1111111111";
                when x"10C3" => data <= "1111111111";
                when x"10C4" => data <= "1111111111";
                when x"10C5" => data <= "1111111111";
                when x"10C6" => data <= "1111111111";
                when x"10C7" => data <= "1111111111";
                when x"10C8" => data <= "1111111111";
                when x"10C9" => data <= "1111111111";
                when x"10CA" => data <= "1111111111";
                when x"10CB" => data <= "1111111111";
                when x"10CC" => data <= "1111111111";
                when x"10CD" => data <= "1111111111";
                when x"10CE" => data <= "0000100100";
                when x"10CF" => data <= "1111111111";
                when x"10D0" => data <= "0010101111";
                when x"10D1" => data <= "1111111111";
                when x"10D2" => data <= "1111111111";
                when x"10D3" => data <= "1111111111";
                when x"10D4" => data <= "1111111111";
                when x"10D5" => data <= "1111111111";
                when x"10D6" => data <= "1111111111";
                when x"10D7" => data <= "1111111111";
                when x"10D8" => data <= "1111111111";
                when x"10D9" => data <= "1111111111";
                when x"10DA" => data <= "1111111111";
                when x"10DB" => data <= "1111111111";
                when x"10DC" => data <= "1111111111";
                when x"10DD" => data <= "1111111111";
                when x"10DE" => data <= "1111111111";
                when x"10DF" => data <= "1111111111";
                when x"10E0" => data <= "1111111111";
                when x"10E1" => data <= "1111111111";
                when x"10E2" => data <= "1111111111";
                when x"10E3" => data <= "1111111111";
                when x"10E4" => data <= "1111111111";
                when x"10E5" => data <= "1111111111";
                when x"10E6" => data <= "1111111111";
                when x"10E7" => data <= "1111111111";
                when x"10E8" => data <= "1111111111";
                when x"10E9" => data <= "1111111111";
                when x"10EA" => data <= "1111111111";
                when x"10EB" => data <= "1111111111";
                when x"10EC" => data <= "1111111111";
                when x"10ED" => data <= "1111111111";
                when x"10EE" => data <= "1111111111";
                when x"10EF" => data <= "1111111111";
                when x"10F0" => data <= "1111111111";
                when x"10F1" => data <= "1111111111";
                when x"10F2" => data <= "1111111111";
                when x"10F3" => data <= "1111111111";
                when x"10F4" => data <= "1111111111";
                when x"10F5" => data <= "1111111111";
                when x"10F6" => data <= "1111111111";
                when x"10F7" => data <= "1111111111";
                when x"10F8" => data <= "1111111111";
                when x"10F9" => data <= "1111111111";
                when x"10FA" => data <= "1111111111";
                when x"10FB" => data <= "1111111111";
                when x"10FC" => data <= "1111111111";
                when x"10FD" => data <= "1111111111";
                when x"10FE" => data <= "1111111111";
                when x"10FF" => data <= "1111111111";
                when x"1100" => data <= "1111111111";
                when x"1101" => data <= "1111111111";
                when x"1102" => data <= "1111111111";
                when x"1103" => data <= "1111111111";
                when x"1104" => data <= "1111111111";
                when x"1105" => data <= "1111111111";
                when x"1106" => data <= "1111111111";
                when x"1107" => data <= "1111111111";
                when x"1108" => data <= "1111111111";
                when x"1109" => data <= "1111111111";
                when x"110A" => data <= "0000100100";
                when x"110B" => data <= "1111111111";
                when x"110C" => data <= "1111111111";
                when x"110D" => data <= "1111111111";
                when x"110E" => data <= "1111111111";
                when x"110F" => data <= "1111111111";
                when x"1110" => data <= "1111111111";
                when x"1111" => data <= "1111111111";
                when x"1112" => data <= "1111111111";
                when x"1113" => data <= "1111111111";
                when x"1114" => data <= "1111111111";
                when x"1115" => data <= "1111111111";
                when x"1116" => data <= "1111111111";
                when x"1117" => data <= "1111111111";
                when x"1118" => data <= "1111111111";
                when x"1119" => data <= "1111111111";
                when x"111A" => data <= "1111111111";
                when x"111B" => data <= "1111111111";
                when x"111C" => data <= "1111111111";
                when x"111D" => data <= "1111111111";
                when x"111E" => data <= "1111111111";
                when x"111F" => data <= "1111111111";
                when x"1120" => data <= "1111111111";
                when x"1121" => data <= "1111111111";
                when x"1122" => data <= "1111111111";
                when x"1123" => data <= "1111111111";
                when x"1124" => data <= "1111111111";
                when x"1125" => data <= "1111111111";
                when x"1126" => data <= "1111111111";
                when x"1127" => data <= "1111111111";
                when x"1128" => data <= "1111111111";
                when x"1129" => data <= "1111111111";
                when x"112A" => data <= "1111111111";
                when x"112B" => data <= "1111111111";
                when x"112C" => data <= "1111111111";
                when x"112D" => data <= "1111111111";
                when x"112E" => data <= "1111111111";
                when x"112F" => data <= "1111111111";
                when x"1130" => data <= "1111111111";
                when x"1131" => data <= "1111111111";
                when x"1132" => data <= "1111111111";
                when x"1133" => data <= "1111111111";
                when x"1134" => data <= "1111111111";
                when x"1135" => data <= "1111111111";
                when x"1136" => data <= "1111111111";
                when x"1137" => data <= "1111111111";
                when x"1138" => data <= "1111111111";
                when x"1139" => data <= "1111111111";
                when x"113A" => data <= "1111111111";
                when x"113B" => data <= "1111111111";
                when x"113C" => data <= "1111111111";
                when x"113D" => data <= "1111111111";
                when x"113E" => data <= "1111111111";
                when x"113F" => data <= "1111111111";
                when x"1140" => data <= "1111111111";
                when x"1141" => data <= "1111111111";
                when x"1142" => data <= "1111111111";
                when x"1143" => data <= "1111111111";
                when x"1144" => data <= "1111111111";
                when x"1145" => data <= "1111111111";
                when x"1146" => data <= "1111111111";
                when x"1147" => data <= "1111111111";
                when x"1148" => data <= "1111111111";
                when x"1149" => data <= "1111111111";
                when x"114A" => data <= "1111111111";
                when x"114B" => data <= "1111111111";
                when x"114C" => data <= "1111111111";
                when x"114D" => data <= "1111111111";
                when x"114E" => data <= "1111111111";
                when x"114F" => data <= "1111111111";
                when x"1150" => data <= "1111111111";
                when x"1151" => data <= "1111111111";
                when x"1152" => data <= "1111111111";
                when x"1153" => data <= "1111111111";
                when x"1154" => data <= "1111111111";
                when x"1155" => data <= "1000001000";
                when x"1156" => data <= "1111111111";
                when x"1157" => data <= "1111111111";
                when x"1158" => data <= "1111111111";
                when x"1159" => data <= "1111111111";
                when x"115A" => data <= "1111111111";
                when x"115B" => data <= "1111111111";
                when x"115C" => data <= "1111111111";
                when x"115D" => data <= "1111111111";
                when x"115E" => data <= "1111111111";
                when x"115F" => data <= "1111111111";
                when x"1160" => data <= "0001111011";
                when x"1161" => data <= "1111111111";
                when x"1162" => data <= "1111111111";
                when x"1163" => data <= "1111111111";
                when x"1164" => data <= "1111111111";
                when x"1165" => data <= "1111111111";
                when x"1166" => data <= "1111111111";
                when x"1167" => data <= "1111111111";
                when x"1168" => data <= "1111111111";
                when x"1169" => data <= "1111111111";
                when x"116A" => data <= "0100000111";
                when x"116B" => data <= "1111111111";
                when x"116C" => data <= "1111111111";
                when x"116D" => data <= "1111111111";
                when x"116E" => data <= "1111111111";
                when x"116F" => data <= "1111111111";
                when x"1170" => data <= "1111111111";
                when x"1171" => data <= "1111111111";
                when x"1172" => data <= "1111111111";
                when x"1173" => data <= "1111111111";
                when x"1174" => data <= "1111111111";
                when x"1175" => data <= "1111111111";
                when x"1176" => data <= "1111111111";
                when x"1177" => data <= "1111111111";
                when x"1178" => data <= "1111111111";
                when x"1179" => data <= "1111111111";
                when x"117A" => data <= "1111111111";
                when x"117B" => data <= "1111111111";
                when x"117C" => data <= "1111111111";
                when x"117D" => data <= "1111111111";
                when x"117E" => data <= "1111111111";
                when x"117F" => data <= "1111111111";
                when x"1180" => data <= "1111111111";
                when x"1181" => data <= "1111111111";
                when x"1182" => data <= "1111111111";
                when x"1183" => data <= "1111111111";
                when x"1184" => data <= "1111111111";
                when x"1185" => data <= "1111111111";
                when x"1186" => data <= "1111111111";
                when x"1187" => data <= "1111111111";
                when x"1188" => data <= "1111111111";
                when x"1189" => data <= "1111111111";
                when x"118A" => data <= "1111111111";
                when x"118B" => data <= "1111111111";
                when x"118C" => data <= "1111111111";
                when x"118D" => data <= "1111111111";
                when x"118E" => data <= "1111111111";
                when x"118F" => data <= "1111111111";
                when x"1190" => data <= "1111111111";
                when x"1191" => data <= "1111111111";
                when x"1192" => data <= "1111111111";
                when x"1193" => data <= "1111111111";
                when x"1194" => data <= "1111111111";
                when x"1195" => data <= "1111111111";
                when x"1196" => data <= "1111111111";
                when x"1197" => data <= "1111111111";
                when x"1198" => data <= "1111111111";
                when x"1199" => data <= "1111111111";
                when x"119A" => data <= "1111111111";
                when x"119B" => data <= "1111111111";
                when x"119C" => data <= "1111111111";
                when x"119D" => data <= "1111111111";
                when x"119E" => data <= "1111111111";
                when x"119F" => data <= "1111111111";
                when x"11A0" => data <= "1111111111";
                when x"11A1" => data <= "1111111111";
                when x"11A2" => data <= "1111111111";
                when x"11A3" => data <= "1111111111";
                when x"11A4" => data <= "1111111111";
                when x"11A5" => data <= "1111111111";
                when x"11A6" => data <= "1111111111";
                when x"11A7" => data <= "1111111111";
                when x"11A8" => data <= "1111111111";
                when x"11A9" => data <= "1111111111";
                when x"11AA" => data <= "1111111111";
                when x"11AB" => data <= "1111111111";
                when x"11AC" => data <= "1111111111";
                when x"11AD" => data <= "1111111111";
                when x"11AE" => data <= "1111111111";
                when x"11AF" => data <= "1111111111";
                when x"11B0" => data <= "1111111111";
                when x"11B1" => data <= "1111111111";
                when x"11B2" => data <= "1111111111";
                when x"11B3" => data <= "1111111111";
                when x"11B4" => data <= "1111111111";
                when x"11B5" => data <= "1111111111";
                when x"11B6" => data <= "1111111111";
                when x"11B7" => data <= "1111111111";
                when x"11B8" => data <= "1111111111";
                when x"11B9" => data <= "1111111111";
                when x"11BA" => data <= "1111111111";
                when x"11BB" => data <= "1111111111";
                when x"11BC" => data <= "1111111111";
                when x"11BD" => data <= "1111111111";
                when x"11BE" => data <= "1111111111";
                when x"11BF" => data <= "1111111111";
                when x"11C0" => data <= "1111111111";
                when x"11C1" => data <= "1111111111";
                when x"11C2" => data <= "1111111111";
                when x"11C3" => data <= "1111111111";
                when x"11C4" => data <= "1111111111";
                when x"11C5" => data <= "1111111111";
                when x"11C6" => data <= "1111111111";
                when x"11C7" => data <= "1111111111";
                when x"11C8" => data <= "1111111111";
                when x"11C9" => data <= "1111111111";
                when x"11CA" => data <= "1111111111";
                when x"11CB" => data <= "1111111111";
                when x"11CC" => data <= "1111111111";
                when x"11CD" => data <= "1111111111";
                when x"11CE" => data <= "1111111111";
                when x"11CF" => data <= "1111111111";
                when x"11D0" => data <= "1111111111";
                when x"11D1" => data <= "1111111111";
                when x"11D2" => data <= "1111111111";
                when x"11D3" => data <= "1111111111";
                when x"11D4" => data <= "1111111111";
                when x"11D5" => data <= "1111111111";
                when x"11D6" => data <= "1111111111";
                when x"11D7" => data <= "1111111111";
                when x"11D8" => data <= "1111111111";
                when x"11D9" => data <= "1111111111";
                when x"11DA" => data <= "1111111111";
                when x"11DB" => data <= "1111111111";
                when x"11DC" => data <= "1111111111";
                when x"11DD" => data <= "1111111111";
                when x"11DE" => data <= "1111111111";
                when x"11DF" => data <= "1111111111";
                when x"11E0" => data <= "1111111111";
                when x"11E1" => data <= "1111111111";
                when x"11E2" => data <= "1111111111";
                when x"11E3" => data <= "1111111111";
                when x"11E4" => data <= "1111111111";
                when x"11E5" => data <= "1111111111";
                when x"11E6" => data <= "1111111111";
                when x"11E7" => data <= "1111111111";
                when x"11E8" => data <= "1111111111";
                when x"11E9" => data <= "1111111111";
                when x"11EA" => data <= "1111111111";
                when x"11EB" => data <= "1111111111";
                when x"11EC" => data <= "1111111111";
                when x"11ED" => data <= "1111111111";
                when x"11EE" => data <= "1111111111";
                when x"11EF" => data <= "1111111111";
                when x"11F0" => data <= "1111111111";
                when x"11F1" => data <= "1111111111";
                when x"11F2" => data <= "1111111111";
                when x"11F3" => data <= "1111111111";
                when x"11F4" => data <= "1111111111";
                when x"11F5" => data <= "1111111111";
                when x"11F6" => data <= "1111111111";
                when x"11F7" => data <= "1111111111";
                when x"11F8" => data <= "1111111111";
                when x"11F9" => data <= "1111111111";
                when x"11FA" => data <= "1111111111";
                when x"11FB" => data <= "1111111111";
                when x"11FC" => data <= "1111111111";
                when x"11FD" => data <= "1111111111";
                when x"11FE" => data <= "1111111111";
                when x"11FF" => data <= "1111111111";
                when x"1200" => data <= "1111111111";
                when x"1201" => data <= "1111111111";
                when x"1202" => data <= "1111111111";
                when x"1203" => data <= "1111111111";
                when x"1204" => data <= "1111111111";
                when x"1205" => data <= "1111111111";
                when x"1206" => data <= "1111111111";
                when x"1207" => data <= "1111111111";
                when x"1208" => data <= "1111111111";
                when x"1209" => data <= "1111111111";
                when x"120A" => data <= "1111111111";
                when x"120B" => data <= "1111111111";
                when x"120C" => data <= "1111111111";
                when x"120D" => data <= "1111111111";
                when x"120E" => data <= "1111111111";
                when x"120F" => data <= "1111111111";
                when x"1210" => data <= "1111111111";
                when x"1211" => data <= "1111111111";
                when x"1212" => data <= "1000111101";
                when x"1213" => data <= "1111111111";
                when x"1214" => data <= "1111111111";
                when x"1215" => data <= "1111111111";
                when x"1216" => data <= "1111111111";
                when x"1217" => data <= "1111111111";
                when x"1218" => data <= "1111111111";
                when x"1219" => data <= "1111111111";
                when x"121A" => data <= "1111111111";
                when x"121B" => data <= "1111111111";
                when x"121C" => data <= "1111111111";
                when x"121D" => data <= "1111111111";
                when x"121E" => data <= "1111111111";
                when x"121F" => data <= "1111111111";
                when x"1220" => data <= "1111111111";
                when x"1221" => data <= "1111111111";
                when x"1222" => data <= "1111111111";
                when x"1223" => data <= "1111111111";
                when x"1224" => data <= "1111111111";
                when x"1225" => data <= "1111111111";
                when x"1226" => data <= "1111111111";
                when x"1227" => data <= "1111111111";
                when x"1228" => data <= "1111111111";
                when x"1229" => data <= "1111111111";
                when x"122A" => data <= "1111111111";
                when x"122B" => data <= "1111111111";
                when x"122C" => data <= "1111111111";
                when x"122D" => data <= "1111111111";
                when x"122E" => data <= "1111111111";
                when x"122F" => data <= "1111111111";
                when x"1230" => data <= "1111111111";
                when x"1231" => data <= "1111111111";
                when x"1232" => data <= "1111111111";
                when x"1233" => data <= "1111111111";
                when x"1234" => data <= "1111111111";
                when x"1235" => data <= "1111111111";
                when x"1236" => data <= "1111111111";
                when x"1237" => data <= "1111111111";
                when x"1238" => data <= "1111111111";
                when x"1239" => data <= "1111111111";
                when x"123A" => data <= "1111111111";
                when x"123B" => data <= "1111111111";
                when x"123C" => data <= "1111111111";
                when x"123D" => data <= "1111111111";
                when x"123E" => data <= "1111111111";
                when x"123F" => data <= "1111111111";
                when x"1240" => data <= "1111111111";
                when x"1241" => data <= "1111111111";
                when x"1242" => data <= "1111111111";
                when x"1243" => data <= "1111111111";
                when x"1244" => data <= "1111111111";
                when x"1245" => data <= "1111111111";
                when x"1246" => data <= "1111111111";
                when x"1247" => data <= "1111111111";
                when x"1248" => data <= "1111111111";
                when x"1249" => data <= "1111111111";
                when x"124A" => data <= "1111111111";
                when x"124B" => data <= "1111111111";
                when x"124C" => data <= "1111111111";
                when x"124D" => data <= "1111111111";
                when x"124E" => data <= "1111111111";
                when x"124F" => data <= "1111111111";
                when x"1250" => data <= "1111111111";
                when x"1251" => data <= "1111111111";
                when x"1252" => data <= "1111111111";
                when x"1253" => data <= "1000001000";
                when x"1254" => data <= "1111111111";
                when x"1255" => data <= "1111111111";
                when x"1256" => data <= "1111111111";
                when x"1257" => data <= "1111111111";
                when x"1258" => data <= "1111111111";
                when x"1259" => data <= "1111111111";
                when x"125A" => data <= "1111111111";
                when x"125B" => data <= "1111111111";
                when x"125C" => data <= "1111111111";
                when x"125D" => data <= "1111111111";
                when x"125E" => data <= "1111111111";
                when x"125F" => data <= "1111111111";
                when x"1260" => data <= "1111111111";
                when x"1261" => data <= "1111111111";
                when x"1262" => data <= "1111111111";
                when x"1263" => data <= "1111111111";
                when x"1264" => data <= "1111111111";
                when x"1265" => data <= "1111111111";
                when x"1266" => data <= "0010101111";
                when x"1267" => data <= "1111111111";
                when x"1268" => data <= "1111111111";
                when x"1269" => data <= "1111111111";
                when x"126A" => data <= "1111111111";
                when x"126B" => data <= "1111111111";
                when x"126C" => data <= "1111111111";
                when x"126D" => data <= "1111111111";
                when x"126E" => data <= "1111111111";
                when x"126F" => data <= "1111111111";
                when x"1270" => data <= "1111111111";
                when x"1271" => data <= "1111111111";
                when x"1272" => data <= "1111111111";
                when x"1273" => data <= "1111111111";
                when x"1274" => data <= "1111111111";
                when x"1275" => data <= "1111111111";
                when x"1276" => data <= "1111111111";
                when x"1277" => data <= "1111111111";
                when x"1278" => data <= "1111111111";
                when x"1279" => data <= "1111111111";
                when x"127A" => data <= "1111111111";
                when x"127B" => data <= "1111111111";
                when x"127C" => data <= "1111111111";
                when x"127D" => data <= "1111111111";
                when x"127E" => data <= "1111111111";
                when x"127F" => data <= "1111111111";
                when x"1280" => data <= "1111111111";
                when x"1281" => data <= "1111111111";
                when x"1282" => data <= "1111111111";
                when x"1283" => data <= "1111111111";
                when x"1284" => data <= "1111111111";
                when x"1285" => data <= "1111111111";
                when x"1286" => data <= "1111111111";
                when x"1287" => data <= "1111111111";
                when x"1288" => data <= "1111111111";
                when x"1289" => data <= "1111111111";
                when x"128A" => data <= "1111111111";
                when x"128B" => data <= "1111111111";
                when x"128C" => data <= "1111111111";
                when x"128D" => data <= "1111111111";
                when x"128E" => data <= "1111111111";
                when x"128F" => data <= "1111111111";
                when x"1290" => data <= "1111111111";
                when x"1291" => data <= "1111111111";
                when x"1292" => data <= "1111111111";
                when x"1293" => data <= "1111111111";
                when x"1294" => data <= "1111111111";
                when x"1295" => data <= "1111111111";
                when x"1296" => data <= "1111111111";
                when x"1297" => data <= "1111111111";
                when x"1298" => data <= "1111111111";
                when x"1299" => data <= "1111111111";
                when x"129A" => data <= "1111111111";
                when x"129B" => data <= "1111111111";
                when x"129C" => data <= "1111111111";
                when x"129D" => data <= "1111111111";
                when x"129E" => data <= "1111111111";
                when x"129F" => data <= "1111111111";
                when x"12A0" => data <= "1111111111";
                when x"12A1" => data <= "1111111111";
                when x"12A2" => data <= "1111111111";
                when x"12A3" => data <= "1111111111";
                when x"12A4" => data <= "1111111111";
                when x"12A5" => data <= "1111111111";
                when x"12A6" => data <= "1111111111";
                when x"12A7" => data <= "1111111111";
                when x"12A8" => data <= "1111111111";
                when x"12A9" => data <= "1111111111";
                when x"12AA" => data <= "1111111111";
                when x"12AB" => data <= "1111111111";
                when x"12AC" => data <= "0000100100";
                when x"12AD" => data <= "1111111111";
                when x"12AE" => data <= "1111111111";
                when x"12AF" => data <= "1111111111";
                when x"12B0" => data <= "1111111111";
                when x"12B1" => data <= "1111111111";
                when x"12B2" => data <= "1111111111";
                when x"12B3" => data <= "1111111111";
                when x"12B4" => data <= "1111111111";
                when x"12B5" => data <= "1111111111";
                when x"12B6" => data <= "1111111111";
                when x"12B7" => data <= "1111111111";
                when x"12B8" => data <= "1111111111";
                when x"12B9" => data <= "1111111111";
                when x"12BA" => data <= "1111111111";
                when x"12BB" => data <= "1111111111";
                when x"12BC" => data <= "1111111111";
                when x"12BD" => data <= "1111111111";
                when x"12BE" => data <= "1111111111";
                when x"12BF" => data <= "1111111111";
                when x"12C0" => data <= "1111111111";
                when x"12C1" => data <= "1111111111";
                when x"12C2" => data <= "1111111111";
                when x"12C3" => data <= "1111111111";
                when x"12C4" => data <= "1111111111";
                when x"12C5" => data <= "1111111111";
                when x"12C6" => data <= "1111111111";
                when x"12C7" => data <= "1111111111";
                when x"12C8" => data <= "1111111111";
                when x"12C9" => data <= "1111111111";
                when x"12CA" => data <= "1111111111";
                when x"12CB" => data <= "1111111111";
                when x"12CC" => data <= "1111111111";
                when x"12CD" => data <= "1111111111";
                when x"12CE" => data <= "1111111111";
                when x"12CF" => data <= "1111111111";
                when x"12D0" => data <= "1111111111";
                when x"12D1" => data <= "1111111111";
                when x"12D2" => data <= "1111111111";
                when x"12D3" => data <= "1111111111";
                when x"12D4" => data <= "1111111111";
                when x"12D5" => data <= "1111111111";
                when x"12D6" => data <= "1111111111";
                when x"12D7" => data <= "1111111111";
                when x"12D8" => data <= "1111111111";
                when x"12D9" => data <= "1111111111";
                when x"12DA" => data <= "1111111111";
                when x"12DB" => data <= "1111111111";
                when x"12DC" => data <= "1111111111";
                when x"12DD" => data <= "1111111111";
                when x"12DE" => data <= "1111111111";
                when x"12DF" => data <= "1111111111";
                when x"12E0" => data <= "1111111111";
                when x"12E1" => data <= "1111111111";
                when x"12E2" => data <= "1111111111";
                when x"12E3" => data <= "1111111111";
                when x"12E4" => data <= "1111111111";
                when x"12E5" => data <= "1111111111";
                when x"12E6" => data <= "1111111111";
                when x"12E7" => data <= "1111111111";
                when x"12E8" => data <= "1111111111";
                when x"12E9" => data <= "1011101001";
                when x"12EA" => data <= "1111111111";
                when x"12EB" => data <= "1111111111";
                when x"12EC" => data <= "1111111111";
                when x"12ED" => data <= "1111111111";
                when x"12EE" => data <= "1111111111";
                when x"12EF" => data <= "1111111111";
                when x"12F0" => data <= "1111111111";
                when x"12F1" => data <= "1111111111";
                when x"12F2" => data <= "1111111111";
                when x"12F3" => data <= "1111111111";
                when x"12F4" => data <= "1111111111";
                when x"12F5" => data <= "1111111111";
                when x"12F6" => data <= "1111111111";
                when x"12F7" => data <= "1111111111";
                when x"12F8" => data <= "1111111111";
                when x"12F9" => data <= "1111111111";
                when x"12FA" => data <= "1111111111";
                when x"12FB" => data <= "1111111111";
                when x"12FC" => data <= "1111111111";
                when x"12FD" => data <= "1111111111";
                when x"12FE" => data <= "1111111111";
                when x"12FF" => data <= "1111111111";
                when x"1300" => data <= "1111111111";
                when x"1301" => data <= "1111111111";
                when x"1302" => data <= "1111111111";
                when x"1303" => data <= "1111111111";
                when x"1304" => data <= "1111111111";
                when x"1305" => data <= "1111111111";
                when x"1306" => data <= "1111111111";
                when x"1307" => data <= "1111111111";
                when x"1308" => data <= "1111111111";
                when x"1309" => data <= "1111111111";
                when x"130A" => data <= "1111111111";
                when x"130B" => data <= "1111111111";
                when x"130C" => data <= "1111111111";
                when x"130D" => data <= "1111111111";
                when x"130E" => data <= "1111111111";
                when x"130F" => data <= "1111111111";
                when x"1310" => data <= "1111111111";
                when x"1311" => data <= "1111111111";
                when x"1312" => data <= "1111111111";
                when x"1313" => data <= "1111111111";
                when x"1314" => data <= "1111111111";
                when x"1315" => data <= "1111111111";
                when x"1316" => data <= "1111111111";
                when x"1317" => data <= "1111111111";
                when x"1318" => data <= "1111111111";
                when x"1319" => data <= "1111111111";
                when x"131A" => data <= "1111111111";
                when x"131B" => data <= "1111111111";
                when x"131C" => data <= "1111111111";
                when x"131D" => data <= "1111111111";
                when x"131E" => data <= "1111111111";
                when x"131F" => data <= "1111111111";
                when x"1320" => data <= "1111111111";
                when x"1321" => data <= "1111111111";
                when x"1322" => data <= "1111111111";
                when x"1323" => data <= "1111111111";
                when x"1324" => data <= "1111111111";
                when x"1325" => data <= "1111111111";
                when x"1326" => data <= "1111111111";
                when x"1327" => data <= "1111111111";
                when x"1328" => data <= "1111111111";
                when x"1329" => data <= "1111111111";
                when x"132A" => data <= "1111111111";
                when x"132B" => data <= "1111111111";
                when x"132C" => data <= "1111111111";
                when x"132D" => data <= "1111111111";
                when x"132E" => data <= "1111111111";
                when x"132F" => data <= "1111111111";
                when x"1330" => data <= "1111111111";
                when x"1331" => data <= "1111111111";
                when x"1332" => data <= "1111111111";
                when x"1333" => data <= "1111111111";
                when x"1334" => data <= "1111111111";
                when x"1335" => data <= "1111111111";
                when x"1336" => data <= "1111111111";
                when x"1337" => data <= "1111111111";
                when x"1338" => data <= "1111111111";
                when x"1339" => data <= "1111111111";
                when x"133A" => data <= "1111111111";
                when x"133B" => data <= "1111111111";
                when x"133C" => data <= "1111111111";
                when x"133D" => data <= "1111111111";
                when x"133E" => data <= "1111111111";
                when x"133F" => data <= "1111111111";
                when x"1340" => data <= "1111111111";
                when x"1341" => data <= "1111111111";
                when x"1342" => data <= "1111111111";
                when x"1343" => data <= "1111111111";
                when x"1344" => data <= "1111111111";
                when x"1345" => data <= "1000001000";
                when x"1346" => data <= "1111111111";
                when x"1347" => data <= "1111111111";
                when x"1348" => data <= "1111111111";
                when x"1349" => data <= "1111111111";
                when x"134A" => data <= "1111111111";
                when x"134B" => data <= "1111111111";
                when x"134C" => data <= "1111111111";
                when x"134D" => data <= "1111111111";
                when x"134E" => data <= "1111111111";
                when x"134F" => data <= "1111111111";
                when x"1350" => data <= "1111111111";
                when x"1351" => data <= "1111111111";
                when x"1352" => data <= "1111111111";
                when x"1353" => data <= "1111111111";
                when x"1354" => data <= "1111111111";
                when x"1355" => data <= "1111111111";
                when x"1356" => data <= "1111111111";
                when x"1357" => data <= "1111111111";
                when x"1358" => data <= "1111111111";
                when x"1359" => data <= "1111111111";
                when x"135A" => data <= "1111111111";
                when x"135B" => data <= "1111111111";
                when x"135C" => data <= "1111111111";
                when x"135D" => data <= "1111111111";
                when x"135E" => data <= "1111111111";
                when x"135F" => data <= "1000001000";
                when x"1360" => data <= "1111111111";
                when x"1361" => data <= "1111111111";
                when x"1362" => data <= "1111111111";
                when x"1363" => data <= "1111111111";
                when x"1364" => data <= "1111111111";
                when x"1365" => data <= "1111111111";
                when x"1366" => data <= "1111111111";
                when x"1367" => data <= "1111111111";
                when x"1368" => data <= "1111111111";
                when x"1369" => data <= "1111111111";
                when x"136A" => data <= "1111111111";
                when x"136B" => data <= "1111111111";
                when x"136C" => data <= "1111111111";
                when x"136D" => data <= "1111111111";
                when x"136E" => data <= "1111111111";
                when x"136F" => data <= "1111111111";
                when x"1370" => data <= "1111111111";
                when x"1371" => data <= "1111111111";
                when x"1372" => data <= "1111111111";
                when x"1373" => data <= "1111111111";
                when x"1374" => data <= "1111111111";
                when x"1375" => data <= "1111111111";
                when x"1376" => data <= "1111111111";
                when x"1377" => data <= "1111111111";
                when x"1378" => data <= "1111111111";
                when x"1379" => data <= "1111111111";
                when x"137A" => data <= "1111111111";
                when x"137B" => data <= "1111111111";
                when x"137C" => data <= "1111111111";
                when x"137D" => data <= "0101101101";
                when x"137E" => data <= "1111111111";
                when x"137F" => data <= "1111111111";
                when x"1380" => data <= "1111111111";
                when x"1381" => data <= "1111111111";
                when x"1382" => data <= "1111111111";
                when x"1383" => data <= "1111111111";
                when x"1384" => data <= "1111111111";
                when x"1385" => data <= "1111111111";
                when x"1386" => data <= "1111111111";
                when x"1387" => data <= "1111111111";
                when x"1388" => data <= "1111111111";
                when x"1389" => data <= "1111111111";
                when x"138A" => data <= "1111111111";
                when x"138B" => data <= "1111111111";
                when x"138C" => data <= "1111111111";
                when x"138D" => data <= "1111111111";
                when x"138E" => data <= "1111111111";
                when x"138F" => data <= "1111111111";
                when x"1390" => data <= "1111111111";
                when x"1391" => data <= "1111111111";
                when x"1392" => data <= "1111111111";
                when x"1393" => data <= "1111111111";
                when x"1394" => data <= "1111111111";
                when x"1395" => data <= "1111111111";
                when x"1396" => data <= "1111111111";
                when x"1397" => data <= "1111111111";
                when x"1398" => data <= "1111111111";
                when x"1399" => data <= "1111111111";
                when x"139A" => data <= "1111111111";
                when x"139B" => data <= "1111111111";
                when x"139C" => data <= "1111111111";
                when x"139D" => data <= "1111111111";
                when x"139E" => data <= "1111111111";
                when x"139F" => data <= "1111111111";
                when x"13A0" => data <= "1111111111";
                when x"13A1" => data <= "1111111111";
                when x"13A2" => data <= "1111111111";
                when x"13A3" => data <= "1111111111";
                when x"13A4" => data <= "1111111111";
                when x"13A5" => data <= "1111111111";
                when x"13A6" => data <= "1111111111";
                when x"13A7" => data <= "1111111111";
                when x"13A8" => data <= "1111111111";
                when x"13A9" => data <= "1111111111";
                when x"13AA" => data <= "1111111111";
                when x"13AB" => data <= "1111111111";
                when x"13AC" => data <= "1111111111";
                when x"13AD" => data <= "1111111111";
                when x"13AE" => data <= "1111111111";
                when x"13AF" => data <= "1111111111";
                when x"13B0" => data <= "1111111111";
                when x"13B1" => data <= "1111111111";
                when x"13B2" => data <= "1111111111";
                when x"13B3" => data <= "1111111111";
                when x"13B4" => data <= "1111111111";
                when x"13B5" => data <= "1111111111";
                when x"13B6" => data <= "1111111111";
                when x"13B7" => data <= "1111111111";
                when x"13B8" => data <= "1111111111";
                when x"13B9" => data <= "1111111111";
                when x"13BA" => data <= "1111111111";
                when x"13BB" => data <= "1111111111";
                when x"13BC" => data <= "1111111111";
                when x"13BD" => data <= "1111111111";
                when x"13BE" => data <= "1111111111";
                when x"13BF" => data <= "1111111111";
                when x"13C0" => data <= "1111111111";
                when x"13C1" => data <= "1111111111";
                when x"13C2" => data <= "1111111111";
                when x"13C3" => data <= "1111111111";
                when x"13C4" => data <= "1111111111";
                when x"13C5" => data <= "1111111111";
                when x"13C6" => data <= "1111111111";
                when x"13C7" => data <= "1111111111";
                when x"13C8" => data <= "1111111111";
                when x"13C9" => data <= "1111111111";
                when x"13CA" => data <= "1111111111";
                when x"13CB" => data <= "1111111111";
                when x"13CC" => data <= "1111111111";
                when x"13CD" => data <= "1111111111";
                when x"13CE" => data <= "1111111111";
                when x"13CF" => data <= "1111111111";
                when x"13D0" => data <= "1000001000";
                when x"13D1" => data <= "1111111111";
                when x"13D2" => data <= "1111111111";
                when x"13D3" => data <= "0001111011";
                when x"13D4" => data <= "1111111111";
                when x"13D5" => data <= "1111111111";
                when x"13D6" => data <= "1111111111";
                when x"13D7" => data <= "1111111111";
                when x"13D8" => data <= "1111111111";
                when x"13D9" => data <= "1111111111";
                when x"13DA" => data <= "1111111111";
                when x"13DB" => data <= "1111111111";
                when x"13DC" => data <= "1111111111";
                when x"13DD" => data <= "1000001000";
                when x"13DE" => data <= "1111111111";
                when x"13DF" => data <= "1111111111";
                when x"13E0" => data <= "1111111111";
                when x"13E1" => data <= "1111111111";
                when x"13E2" => data <= "1111111111";
                when x"13E3" => data <= "1111111111";
                when x"13E4" => data <= "1111111111";
                when x"13E5" => data <= "1111111111";
                when x"13E6" => data <= "1111111111";
                when x"13E7" => data <= "1111111111";
                when x"13E8" => data <= "1000001000";
                when x"13E9" => data <= "1111111111";
                when x"13EA" => data <= "1111111111";
                when x"13EB" => data <= "1111111111";
                when x"13EC" => data <= "1111111111";
                when x"13ED" => data <= "1111111111";
                when x"13EE" => data <= "1111111111";
                when x"13EF" => data <= "1111111111";
                when x"13F0" => data <= "1111111111";
                when x"13F1" => data <= "1111111111";
                when x"13F2" => data <= "1111111111";
                when x"13F3" => data <= "1111111111";
                when x"13F4" => data <= "1111111111";
                when x"13F5" => data <= "1111111111";
                when x"13F6" => data <= "1111111111";
                when x"13F7" => data <= "1111111111";
                when x"13F8" => data <= "1111111111";
                when x"13F9" => data <= "1111111111";
                when x"13FA" => data <= "1111111111";
                when x"13FB" => data <= "1111111111";
                when x"13FC" => data <= "1111111111";
                when x"13FD" => data <= "1111111111";
                when x"13FE" => data <= "1111111111";
                when x"13FF" => data <= "1111111111";
                when x"1400" => data <= "1111111111";
                when x"1401" => data <= "1111111111";
                when x"1402" => data <= "1111111111";
                when x"1403" => data <= "1111111111";
                when x"1404" => data <= "1111111111";
                when x"1405" => data <= "1111111111";
                when x"1406" => data <= "1111111111";
                when x"1407" => data <= "1111111111";
                when x"1408" => data <= "1111111111";
                when x"1409" => data <= "1111111111";
                when x"140A" => data <= "1111111111";
                when x"140B" => data <= "1111111111";
                when x"140C" => data <= "1111111111";
                when x"140D" => data <= "1111111111";
                when x"140E" => data <= "1111111111";
                when x"140F" => data <= "1111111111";
                when x"1410" => data <= "1111111111";
                when x"1411" => data <= "1111111111";
                when x"1412" => data <= "1111111111";
                when x"1413" => data <= "1111111111";
                when x"1414" => data <= "1111111111";
                when x"1415" => data <= "1111111111";
                when x"1416" => data <= "1111111111";
                when x"1417" => data <= "1111111111";
                when x"1418" => data <= "1111111111";
                when x"1419" => data <= "1111111111";
                when x"141A" => data <= "1111111111";
                when x"141B" => data <= "1111111111";
                when x"141C" => data <= "1111111111";
                when x"141D" => data <= "1111111111";
                when x"141E" => data <= "1111111111";
                when x"141F" => data <= "1111111111";
                when x"1420" => data <= "1111111111";
                when x"1421" => data <= "1111111111";
                when x"1422" => data <= "1111111111";
                when x"1423" => data <= "1111111111";
                when x"1424" => data <= "1111111111";
                when x"1425" => data <= "1111111111";
                when x"1426" => data <= "1111111111";
                when x"1427" => data <= "1111111111";
                when x"1428" => data <= "1111111111";
                when x"1429" => data <= "1111111111";
                when x"142A" => data <= "1111111111";
                when x"142B" => data <= "1111111111";
                when x"142C" => data <= "1111111111";
                when x"142D" => data <= "1111111111";
                when x"142E" => data <= "1111111111";
                when x"142F" => data <= "1111111111";
                when x"1430" => data <= "1111111111";
                when x"1431" => data <= "1111111111";
                when x"1432" => data <= "1111111111";
                when x"1433" => data <= "1111111111";
                when x"1434" => data <= "1111111111";
                when x"1435" => data <= "1111111111";
                when x"1436" => data <= "1111111111";
                when x"1437" => data <= "1111111111";
                when x"1438" => data <= "1111111111";
                when x"1439" => data <= "1111111111";
                when x"143A" => data <= "1111111111";
                when x"143B" => data <= "1111111111";
                when x"143C" => data <= "1111111111";
                when x"143D" => data <= "1111111111";
                when x"143E" => data <= "1111111111";
                when x"143F" => data <= "1111111111";
                when x"1440" => data <= "1111111111";
                when x"1441" => data <= "1111111111";
                when x"1442" => data <= "1111111111";
                when x"1443" => data <= "1111111111";
                when x"1444" => data <= "1111111111";
                when x"1445" => data <= "1111111111";
                when x"1446" => data <= "1111111111";
                when x"1447" => data <= "1111111111";
                when x"1448" => data <= "1111111111";
                when x"1449" => data <= "1111111111";
                when x"144A" => data <= "1111111111";
                when x"144B" => data <= "1111111111";
                when x"144C" => data <= "1111111111";
                when x"144D" => data <= "1111111111";
                when x"144E" => data <= "1111111111";
                when x"144F" => data <= "1111111111";
                when x"1450" => data <= "1111111111";
                when x"1451" => data <= "1111111111";
                when x"1452" => data <= "1111111111";
                when x"1453" => data <= "1111111111";
                when x"1454" => data <= "1111111111";
                when x"1455" => data <= "1111111111";
                when x"1456" => data <= "1111111111";
                when x"1457" => data <= "1111111111";
                when x"1458" => data <= "1111111111";
                when x"1459" => data <= "1111111111";
                when x"145A" => data <= "1111111111";
                when x"145B" => data <= "1111111111";
                when x"145C" => data <= "1111111111";
                when x"145D" => data <= "1111111111";
                when x"145E" => data <= "1111111111";
                when x"145F" => data <= "1111111111";
                when x"1460" => data <= "1111111111";
                when x"1461" => data <= "1111111111";
                when x"1462" => data <= "1111111111";
                when x"1463" => data <= "1111111111";
                when x"1464" => data <= "1111111111";
                when x"1465" => data <= "1111111111";
                when x"1466" => data <= "1111111111";
                when x"1467" => data <= "1111111111";
                when x"1468" => data <= "1111111111";
                when x"1469" => data <= "0101101101";
                when x"146A" => data <= "1111111111";
                when x"146B" => data <= "1111111111";
                when x"146C" => data <= "1111111111";
                when x"146D" => data <= "1111111111";
                when x"146E" => data <= "1111111111";
                when x"146F" => data <= "1111111111";
                when x"1470" => data <= "1111111111";
                when x"1471" => data <= "1111111111";
                when x"1472" => data <= "1111111111";
                when x"1473" => data <= "1111111111";
                when x"1474" => data <= "1111111111";
                when x"1475" => data <= "1111111111";
                when x"1476" => data <= "1111111111";
                when x"1477" => data <= "1111111111";
                when x"1478" => data <= "1111111111";
                when x"1479" => data <= "1111111111";
                when x"147A" => data <= "1111111111";
                when x"147B" => data <= "1111111111";
                when x"147C" => data <= "1111111111";
                when x"147D" => data <= "1111111111";
                when x"147E" => data <= "1111111111";
                when x"147F" => data <= "1111111111";
                when x"1480" => data <= "1111111111";
                when x"1481" => data <= "1111111111";
                when x"1482" => data <= "1111111111";
                when x"1483" => data <= "1111111111";
                when x"1484" => data <= "1111111111";
                when x"1485" => data <= "1111111111";
                when x"1486" => data <= "1111111111";
                when x"1487" => data <= "1111111111";
                when x"1488" => data <= "1111111111";
                when x"1489" => data <= "1111111111";
                when x"148A" => data <= "1111111111";
                when x"148B" => data <= "1111111111";
                when x"148C" => data <= "1111111111";
                when x"148D" => data <= "1111111111";
                when x"148E" => data <= "1111111111";
                when x"148F" => data <= "1111111111";
                when x"1490" => data <= "1111111111";
                when x"1491" => data <= "1111111111";
                when x"1492" => data <= "1111111111";
                when x"1493" => data <= "1111111111";
                when x"1494" => data <= "1111111111";
                when x"1495" => data <= "1111111111";
                when x"1496" => data <= "1111111111";
                when x"1497" => data <= "1111111111";
                when x"1498" => data <= "1111111111";
                when x"1499" => data <= "1111111111";
                when x"149A" => data <= "1111111111";
                when x"149B" => data <= "1111111111";
                when x"149C" => data <= "1111111111";
                when x"149D" => data <= "1111111111";
                when x"149E" => data <= "1111111111";
                when x"149F" => data <= "1111111111";
                when x"14A0" => data <= "1111111111";
                when x"14A1" => data <= "1111111111";
                when x"14A2" => data <= "1111111111";
                when x"14A3" => data <= "1111111111";
                when x"14A4" => data <= "1111111111";
                when x"14A5" => data <= "1111111111";
                when x"14A6" => data <= "1111111111";
                when x"14A7" => data <= "1111111111";
                when x"14A8" => data <= "1111111111";
                when x"14A9" => data <= "1111111111";
                when x"14AA" => data <= "1111111111";
                when x"14AB" => data <= "1111111111";
                when x"14AC" => data <= "1111111111";
                when x"14AD" => data <= "1111111111";
                when x"14AE" => data <= "1111111111";
                when x"14AF" => data <= "1111111111";
                when x"14B0" => data <= "1111111111";
                when x"14B1" => data <= "1111111111";
                when x"14B2" => data <= "1111111111";
                when x"14B3" => data <= "1111111111";
                when x"14B4" => data <= "1111111111";
                when x"14B5" => data <= "1111111111";
                when x"14B6" => data <= "1111111111";
                when x"14B7" => data <= "1111111111";
                when x"14B8" => data <= "1111111111";
                when x"14B9" => data <= "1111111111";
                when x"14BA" => data <= "1111111111";
                when x"14BB" => data <= "1111111111";
                when x"14BC" => data <= "1111111111";
                when x"14BD" => data <= "1111111111";
                when x"14BE" => data <= "1111111111";
                when x"14BF" => data <= "1111111111";
                when x"14C0" => data <= "1111111111";
                when x"14C1" => data <= "1111111111";
                when x"14C2" => data <= "1111111111";
                when x"14C3" => data <= "1111111111";
                when x"14C4" => data <= "1111111111";
                when x"14C5" => data <= "1111111111";
                when x"14C6" => data <= "1111111111";
                when x"14C7" => data <= "1111111111";
                when x"14C8" => data <= "1111111111";
                when x"14C9" => data <= "1111111111";
                when x"14CA" => data <= "1111111111";
                when x"14CB" => data <= "1111111111";
                when x"14CC" => data <= "1111111111";
                when x"14CD" => data <= "1111111111";
                when x"14CE" => data <= "1111111111";
                when x"14CF" => data <= "1111111111";
                when x"14D0" => data <= "1111111111";
                when x"14D1" => data <= "1111111111";
                when x"14D2" => data <= "1111111111";
                when x"14D3" => data <= "1111111111";
                when x"14D4" => data <= "1111111111";
                when x"14D5" => data <= "1111111111";
                when x"14D6" => data <= "1111111111";
                when x"14D7" => data <= "1111111111";
                when x"14D8" => data <= "1111111111";
                when x"14D9" => data <= "1111111111";
                when x"14DA" => data <= "1111111111";
                when x"14DB" => data <= "1111111111";
                when x"14DC" => data <= "1111111111";
                when x"14DD" => data <= "1111111111";
                when x"14DE" => data <= "1111111111";
                when x"14DF" => data <= "1111111111";
                when x"14E0" => data <= "1111111111";
                when x"14E1" => data <= "1111111111";
                when x"14E2" => data <= "1111111111";
                when x"14E3" => data <= "1111111111";
                when x"14E4" => data <= "1111111111";
                when x"14E5" => data <= "1111111111";
                when x"14E6" => data <= "1111111111";
                when x"14E7" => data <= "1111111111";
                when x"14E8" => data <= "1111111111";
                when x"14E9" => data <= "1111111111";
                when x"14EA" => data <= "1111111111";
                when x"14EB" => data <= "1111111111";
                when x"14EC" => data <= "1111111111";
                when x"14ED" => data <= "1111111111";
                when x"14EE" => data <= "1111111111";
                when x"14EF" => data <= "1111111111";
                when x"14F0" => data <= "1111111111";
                when x"14F1" => data <= "1111111111";
                when x"14F2" => data <= "1111111111";
                when x"14F3" => data <= "1111111111";
                when x"14F4" => data <= "1111111111";
                when x"14F5" => data <= "1111111111";
                when x"14F6" => data <= "1111111111";
                when x"14F7" => data <= "1111111111";
                when x"14F8" => data <= "1111111111";
                when x"14F9" => data <= "1111111111";
                when x"14FA" => data <= "1111111111";
                when x"14FB" => data <= "1111111111";
                when x"14FC" => data <= "1111111111";
                when x"14FD" => data <= "1111111111";
                when x"14FE" => data <= "1111111111";
                when x"14FF" => data <= "1111111111";
                when x"1500" => data <= "1111111111";
                when x"1501" => data <= "1111111111";
                when x"1502" => data <= "1111111111";
                when x"1503" => data <= "1111111111";
                when x"1504" => data <= "1111111111";
                when x"1505" => data <= "1111111111";
                when x"1506" => data <= "1111111111";
                when x"1507" => data <= "1111111111";
                when x"1508" => data <= "1111111111";
                when x"1509" => data <= "1111111111";
                when x"150A" => data <= "1111111111";
                when x"150B" => data <= "1111111111";
                when x"150C" => data <= "1111111111";
                when x"150D" => data <= "1111111111";
                when x"150E" => data <= "1111111111";
                when x"150F" => data <= "1111111111";
                when x"1510" => data <= "1111111111";
                when x"1511" => data <= "1111111111";
                when x"1512" => data <= "1111111111";
                when x"1513" => data <= "1111111111";
                when x"1514" => data <= "1111111111";
                when x"1515" => data <= "1111111111";
                when x"1516" => data <= "1111111111";
                when x"1517" => data <= "1111111111";
                when x"1518" => data <= "1111111111";
                when x"1519" => data <= "1111111111";
                when x"151A" => data <= "1111111111";
                when x"151B" => data <= "1111111111";
                when x"151C" => data <= "1111111111";
                when x"151D" => data <= "1111111111";
                when x"151E" => data <= "1111111111";
                when x"151F" => data <= "1111111111";
                when x"1520" => data <= "1111111111";
                when x"1521" => data <= "1111111111";
                when x"1522" => data <= "1111111111";
                when x"1523" => data <= "1111111111";
                when x"1524" => data <= "0101011000";
                when x"1525" => data <= "1111111111";
                when x"1526" => data <= "1111111111";
                when x"1527" => data <= "1111111111";
                when x"1528" => data <= "1111111111";
                when x"1529" => data <= "1111111111";
                when x"152A" => data <= "1111111111";
                when x"152B" => data <= "1111111111";
                when x"152C" => data <= "1111111111";
                when x"152D" => data <= "1111111111";
                when x"152E" => data <= "1111111111";
                when x"152F" => data <= "1111111111";
                when x"1530" => data <= "1111111111";
                when x"1531" => data <= "1111111111";
                when x"1532" => data <= "1111111111";
                when x"1533" => data <= "1111111111";
                when x"1534" => data <= "1111111111";
                when x"1535" => data <= "1111111111";
                when x"1536" => data <= "1111111111";
                when x"1537" => data <= "1111111111";
                when x"1538" => data <= "1111111111";
                when x"1539" => data <= "1111111111";
                when x"153A" => data <= "1111111111";
                when x"153B" => data <= "1111111111";
                when x"153C" => data <= "1111111111";
                when x"153D" => data <= "1111111111";
                when x"153E" => data <= "1111111111";
                when x"153F" => data <= "1111111111";
                when x"1540" => data <= "1111111111";
                when x"1541" => data <= "1111111111";
                when x"1542" => data <= "1111111111";
                when x"1543" => data <= "1111111111";
                when x"1544" => data <= "1111111111";
                when x"1545" => data <= "1111111111";
                when x"1546" => data <= "1111111111";
                when x"1547" => data <= "1111111111";
                when x"1548" => data <= "1111111111";
                when x"1549" => data <= "1111111111";
                when x"154A" => data <= "1111111111";
                when x"154B" => data <= "1111111111";
                when x"154C" => data <= "1111111111";
                when x"154D" => data <= "1111111111";
                when x"154E" => data <= "1111111111";
                when x"154F" => data <= "1111111111";
                when x"1550" => data <= "1111111111";
                when x"1551" => data <= "1111111111";
                when x"1552" => data <= "1111111111";
                when x"1553" => data <= "1111111111";
                when x"1554" => data <= "1111111111";
                when x"1555" => data <= "1111111111";
                when x"1556" => data <= "1111111111";
                when x"1557" => data <= "1111111111";
                when x"1558" => data <= "1111111111";
                when x"1559" => data <= "1111111111";
                when x"155A" => data <= "1111111111";
                when x"155B" => data <= "1111111111";
                when x"155C" => data <= "1111111111";
                when x"155D" => data <= "1111111111";
                when x"155E" => data <= "1000111101";
                when x"155F" => data <= "1111111111";
                when x"1560" => data <= "1111111111";
                when x"1561" => data <= "1111111111";
                when x"1562" => data <= "1111111111";
                when x"1563" => data <= "1111111111";
                when x"1564" => data <= "1111111111";
                when x"1565" => data <= "1111111111";
                when x"1566" => data <= "1111111111";
                when x"1567" => data <= "1111111111";
                when x"1568" => data <= "1111111111";
                when x"1569" => data <= "1111111111";
                when x"156A" => data <= "1111111111";
                when x"156B" => data <= "1111111111";
                when x"156C" => data <= "1111111111";
                when x"156D" => data <= "1111111111";
                when x"156E" => data <= "1111111111";
                when x"156F" => data <= "1111111111";
                when x"1570" => data <= "1111111111";
                when x"1571" => data <= "1111111111";
                when x"1572" => data <= "1111111111";
                when x"1573" => data <= "1111111111";
                when x"1574" => data <= "1111111111";
                when x"1575" => data <= "1111111111";
                when x"1576" => data <= "1111111111";
                when x"1577" => data <= "1111111111";
                when x"1578" => data <= "1111111111";
                when x"1579" => data <= "1111111111";
                when x"157A" => data <= "1111111111";
                when x"157B" => data <= "1111111111";
                when x"157C" => data <= "1111111111";
                when x"157D" => data <= "1111111111";
                when x"157E" => data <= "1111111111";
                when x"157F" => data <= "1111111111";
                when x"1580" => data <= "1111111111";
                when x"1581" => data <= "1111111111";
                when x"1582" => data <= "1111111111";
                when x"1583" => data <= "1111111111";
                when x"1584" => data <= "1111111111";
                when x"1585" => data <= "1111111111";
                when x"1586" => data <= "1111111111";
                when x"1587" => data <= "1111111111";
                when x"1588" => data <= "1111111111";
                when x"1589" => data <= "1111111111";
                when x"158A" => data <= "1111111111";
                when x"158B" => data <= "1111111111";
                when x"158C" => data <= "1111111111";
                when x"158D" => data <= "1111111111";
                when x"158E" => data <= "1111111111";
                when x"158F" => data <= "1111111111";
                when x"1590" => data <= "1111111111";
                when x"1591" => data <= "1111111111";
                when x"1592" => data <= "1111111111";
                when x"1593" => data <= "1111111111";
                when x"1594" => data <= "1111111111";
                when x"1595" => data <= "1111111111";
                when x"1596" => data <= "1111111111";
                when x"1597" => data <= "1111111111";
                when x"1598" => data <= "1111111111";
                when x"1599" => data <= "1111111111";
                when x"159A" => data <= "1111111111";
                when x"159B" => data <= "1111111111";
                when x"159C" => data <= "1111111111";
                when x"159D" => data <= "1111111111";
                when x"159E" => data <= "1111111111";
                when x"159F" => data <= "1111111111";
                when x"15A0" => data <= "1111111111";
                when x"15A1" => data <= "1111111111";
                when x"15A2" => data <= "1111111111";
                when x"15A3" => data <= "1111111111";
                when x"15A4" => data <= "1111111111";
                when x"15A5" => data <= "1111111111";
                when x"15A6" => data <= "1111111111";
                when x"15A7" => data <= "1111111111";
                when x"15A8" => data <= "1111111111";
                when x"15A9" => data <= "1111111111";
                when x"15AA" => data <= "1111111111";
                when x"15AB" => data <= "1111111111";
                when x"15AC" => data <= "1111111111";
                when x"15AD" => data <= "1111111111";
                when x"15AE" => data <= "1111111111";
                when x"15AF" => data <= "1111111111";
                when x"15B0" => data <= "1111111111";
                when x"15B1" => data <= "1111111111";
                when x"15B2" => data <= "1111111111";
                when x"15B3" => data <= "1111111111";
                when x"15B4" => data <= "1111111111";
                when x"15B5" => data <= "1111111111";
                when x"15B6" => data <= "1111111111";
                when x"15B7" => data <= "1111111111";
                when x"15B8" => data <= "1111111111";
                when x"15B9" => data <= "1111111111";
                when x"15BA" => data <= "1111111111";
                when x"15BB" => data <= "1111111111";
                when x"15BC" => data <= "1111111111";
                when x"15BD" => data <= "1111111111";
                when x"15BE" => data <= "1111111111";
                when x"15BF" => data <= "1111111111";
                when x"15C0" => data <= "1111111111";
                when x"15C1" => data <= "1111111111";
                when x"15C2" => data <= "1111111111";
                when x"15C3" => data <= "1111111111";
                when x"15C4" => data <= "1111111111";
                when x"15C5" => data <= "1111111111";
                when x"15C6" => data <= "1111111111";
                when x"15C7" => data <= "1111111111";
                when x"15C8" => data <= "1111111111";
                when x"15C9" => data <= "1111111111";
                when x"15CA" => data <= "1111111111";
                when x"15CB" => data <= "1111111111";
                when x"15CC" => data <= "1111111111";
                when x"15CD" => data <= "1111111111";
                when x"15CE" => data <= "1111111111";
                when x"15CF" => data <= "1111111111";
                when x"15D0" => data <= "1111111111";
                when x"15D1" => data <= "1111111111";
                when x"15D2" => data <= "1111111111";
                when x"15D3" => data <= "1111111111";
                when x"15D4" => data <= "1111111111";
                when x"15D5" => data <= "1111111111";
                when x"15D6" => data <= "1111111111";
                when x"15D7" => data <= "1111111111";
                when x"15D8" => data <= "1111111111";
                when x"15D9" => data <= "1111111111";
                when x"15DA" => data <= "1111111111";
                when x"15DB" => data <= "1111111111";
                when x"15DC" => data <= "1111111111";
                when x"15DD" => data <= "1111111111";
                when x"15DE" => data <= "1111111111";
                when x"15DF" => data <= "1111111111";
                when x"15E0" => data <= "1111111111";
                when x"15E1" => data <= "1111111111";
                when x"15E2" => data <= "1111111111";
                when x"15E3" => data <= "1111111111";
                when x"15E4" => data <= "1111111111";
                when x"15E5" => data <= "1111111111";
                when x"15E6" => data <= "1111111111";
                when x"15E7" => data <= "1111111111";
                when x"15E8" => data <= "1111111111";
                when x"15E9" => data <= "1111111111";
                when x"15EA" => data <= "1111111111";
                when x"15EB" => data <= "1111111111";
                when x"15EC" => data <= "1111111111";
                when x"15ED" => data <= "1111111111";
                when x"15EE" => data <= "1111111111";
                when x"15EF" => data <= "1111111111";
                when x"15F0" => data <= "1111111111";
                when x"15F1" => data <= "1111111111";
                when x"15F2" => data <= "1111111111";
                when x"15F3" => data <= "1111111111";
                when x"15F4" => data <= "1111111111";
                when x"15F5" => data <= "1111111111";
                when x"15F6" => data <= "1111111111";
                when x"15F7" => data <= "1111111111";
                when x"15F8" => data <= "1111111111";
                when x"15F9" => data <= "1111111111";
                when x"15FA" => data <= "1111111111";
                when x"15FB" => data <= "1111111111";
                when x"15FC" => data <= "1111111111";
                when x"15FD" => data <= "1111111111";
                when x"15FE" => data <= "1111111111";
                when x"15FF" => data <= "0100000111";
                when x"1600" => data <= "1111111111";
                when x"1601" => data <= "1111111111";
                when x"1602" => data <= "1111111111";
                when x"1603" => data <= "1111111111";
                when x"1604" => data <= "1111111111";
                when x"1605" => data <= "1111111111";
                when x"1606" => data <= "1111111111";
                when x"1607" => data <= "1111111111";
                when x"1608" => data <= "1111111111";
                when x"1609" => data <= "1111111111";
                when x"160A" => data <= "1111111111";
                when x"160B" => data <= "1111111111";
                when x"160C" => data <= "1111111111";
                when x"160D" => data <= "1111111111";
                when x"160E" => data <= "1111111111";
                when x"160F" => data <= "1111111111";
                when x"1610" => data <= "1111111111";
                when x"1611" => data <= "1111111111";
                when x"1612" => data <= "1111111111";
                when x"1613" => data <= "1111111111";
                when x"1614" => data <= "1111111111";
                when x"1615" => data <= "1111111111";
                when x"1616" => data <= "1111111111";
                when x"1617" => data <= "1111111111";
                when x"1618" => data <= "1111111111";
                when x"1619" => data <= "1111111111";
                when x"161A" => data <= "1111111111";
                when x"161B" => data <= "1111111111";
                when x"161C" => data <= "1111111111";
                when x"161D" => data <= "1111111111";
                when x"161E" => data <= "1111111111";
                when x"161F" => data <= "1111111111";
                when x"1620" => data <= "1111111111";
                when x"1621" => data <= "1111111111";
                when x"1622" => data <= "1111111111";
                when x"1623" => data <= "1111111111";
                when x"1624" => data <= "1111111111";
                when x"1625" => data <= "1111111111";
                when x"1626" => data <= "1111111111";
                when x"1627" => data <= "1111111111";
                when x"1628" => data <= "1111111111";
                when x"1629" => data <= "1111111111";
                when x"162A" => data <= "1111111111";
                when x"162B" => data <= "1111111111";
                when x"162C" => data <= "1111111111";
                when x"162D" => data <= "1111111111";
                when x"162E" => data <= "1111111111";
                when x"162F" => data <= "1111111111";
                when x"1630" => data <= "1111111111";
                when x"1631" => data <= "1111111111";
                when x"1632" => data <= "1111111111";
                when x"1633" => data <= "1111111111";
                when x"1634" => data <= "1111111111";
                when x"1635" => data <= "1111111111";
                when x"1636" => data <= "1111111111";
                when x"1637" => data <= "0100010000";
                when x"1638" => data <= "1110000010";
                when x"1639" => data <= "1001000000";
                when x"163A" => data <= "0011010010";
                when x"163B" => data <= "1101010110";
                when x"163C" => data <= "1001000000";
                when x"163D" => data <= "0110101110";
                when x"163E" => data <= "1001000000";
                when x"163F" => data <= "1111011101";
                when x"1640" => data <= "1001000000";
                when x"1641" => data <= "0100100101";
                when x"1642" => data <= "1001000000";
                when x"1643" => data <= "0100100101";
                when x"1644" => data <= "0100100101";
                when x"1645" => data <= "0100100101";
                when x"1646" => data <= "0000000110";
                when x"1647" => data <= "1101010110";
                when x"1648" => data <= "1110110111";
                when x"1649" => data <= "0100100101";
                when x"164A" => data <= "0100100101";
                when x"164B" => data <= "0100010000";
                when x"164C" => data <= "1101010110";
                when x"164D" => data <= "1111101000";
                when x"164E" => data <= "1111011101";
                when x"164F" => data <= "0100100101";
                when x"1650" => data <= "1001000000";
                when x"1651" => data <= "1001000000";
                when x"1652" => data <= "1001110101";
                when x"1653" => data <= "1000011111";
                when x"1654" => data <= "0100100101";
                when x"1655" => data <= "1001000000";
                when x"1656" => data <= "1001000000";
                when x"1657" => data <= "1010100001";
                when x"1658" => data <= "1001000000";
                when x"1659" => data <= "0111000100";
                when x"165A" => data <= "1001000000";
                when x"165B" => data <= "1110000010";
                when x"165C" => data <= "1001000000";
                when x"165D" => data <= "1001110101";
                when x"165E" => data <= "1001000000";
                when x"165F" => data <= "1001000000";
                when x"1660" => data <= "1101010110";
                when x"1661" => data <= "0100100101";
                when x"1662" => data <= "1000101010";
                when x"1663" => data <= "1001000000";
                when x"1664" => data <= "1001000000";
                when x"1665" => data <= "0100100101";
                when x"1666" => data <= "0100010000";
                when x"1667" => data <= "1001000000";
                when x"1668" => data <= "0100100101";
                when x"1669" => data <= "1101010110";
                when x"166A" => data <= "0100010000";
                when x"166B" => data <= "0100010000";
                when x"166C" => data <= "1001000000";
                when x"166D" => data <= "1001000000";
                when x"166E" => data <= "1000101010";
                when x"166F" => data <= "0100100101";
                when x"1670" => data <= "1000000101";
                when x"1671" => data <= "1110011000";
                when x"1672" => data <= "1100010011";
                when x"1673" => data <= "0111101011";
                when x"1674" => data <= "1110011000";
                when x"1675" => data <= "1110011000";
                when x"1676" => data <= "0100111111";
                when x"1677" => data <= "1110101101";
                when x"1678" => data <= "1111110010";
                when x"1679" => data <= "1010001110";
                when x"167A" => data <= "1111110010";
                when x"167B" => data <= "1010111011";
                when x"167C" => data <= "0100001010";
                when x"167D" => data <= "1000110000";
                when x"167E" => data <= "0100111111";
                when x"167F" => data <= "1101111001";
                when x"1680" => data <= "0000101001";
                when x"1681" => data <= "0000101001";
                when x"1682" => data <= "0101010101";
                when x"1683" => data <= "1000000101";
                when x"1684" => data <= "1110101101";
                when x"1685" => data <= "0100111111";
                when x"1686" => data <= "0100001010";
                when x"1687" => data <= "1111000111";
                when x"1688" => data <= "0110000001";
                when x"1689" => data <= "0100111111";
                when x"168A" => data <= "1001011010";
                when x"168B" => data <= "1010111011";
                when x"168C" => data <= "0111011110";
                when x"168D" => data <= "1001011010";
                when x"168E" => data <= "0101010101";
                when x"168F" => data <= "1111110010";
                when x"1690" => data <= "0001000011";
                when x"1691" => data <= "1001101111";
                when x"1692" => data <= "0111011110";
                when x"1693" => data <= "0101010101";
                when x"1694" => data <= "1000000101";
                when x"1695" => data <= "1011100100";
                when x"1696" => data <= "0011001000";
                when x"1697" => data <= "1000000101";
                when x"1698" => data <= "0001110110";
                when x"1699" => data <= "1110101101";
                when x"169A" => data <= "0111011110";
                when x"169B" => data <= "0000101001";
                when x"169C" => data <= "0111101011";
                when x"169D" => data <= "1001100100";
                when x"169E" => data <= "1011011010";
                when x"169F" => data <= "1100011000";
                when x"16A0" => data <= "1011011010";
                when x"16A1" => data <= "0110001010";
                when x"16A2" => data <= "1011101111";
                when x"16A3" => data <= "0110001010";
                when x"16A4" => data <= "0010101001";
                when x"16A5" => data <= "1000111011";
                when x"16A6" => data <= "1011011010";
                when x"16A7" => data <= "0001001000";
                when x"16A8" => data <= "1111001100";
                when x"16A9" => data <= "0111100000";
                when x"16AA" => data <= "0010101001";
                when x"16AB" => data <= "0000100010";
                when x"16AC" => data <= "0110111111";
                when x"16AD" => data <= "1011011010";
                when x"16AE" => data <= "1111111001";
                when x"16AF" => data <= "1011011010";
                when x"16B0" => data <= "0001111101";
                when x"16B1" => data <= "0110001010";
                when x"16B2" => data <= "0000100010";
                when x"16B3" => data <= "0110001010";
                when x"16B4" => data <= "0110111111";
                when x"16B5" => data <= "0110111111";
                when x"16B6" => data <= "0110111111";
                when x"16B7" => data <= "1011101111";
                when x"16B8" => data <= "0110111111";
                when x"16B9" => data <= "1011011010";
                when x"16BA" => data <= "0110111111";
                when x"16BB" => data <= "0110111111";
                when x"16BC" => data <= "0010101001";
                when x"16BD" => data <= "0000100010";
                when x"16BE" => data <= "0110001010";
                when x"16BF" => data <= "0110111111";
                when x"16C0" => data <= "0000010111";
                when x"16C1" => data <= "0110111111";
                when x"16C2" => data <= "1011011010";
                when x"16C3" => data <= "0111010101";
                when x"16C4" => data <= "1011011010";
                when x"16C5" => data <= "1011101111";
                when x"16C6" => data <= "0101011110";
                when x"16C7" => data <= "0110111111";
                when x"16C8" => data <= "0100000001";
                when x"16C9" => data <= "0110111111";
                when x"16CA" => data <= "0111010101";
                when x"16CB" => data <= "1011011010";
                when x"16CC" => data <= "0100000001";
                when x"16CD" => data <= "1010000101";
                when x"16CE" => data <= "0001001000";
                when x"16CF" => data <= "0001001000";
                when x"16D0" => data <= "0110111111";
                when x"16D1" => data <= "0110001010";
                when x"16D2" => data <= "0110001010";
                when x"16D3" => data <= "1101110010";
                when x"16D4" => data <= "0000100010";
                when x"16D5" => data <= "0110111111";
                when x"16D6" => data <= "0010101001";
                when x"16D7" => data <= "0000100010";
                when x"16D8" => data <= "1011011010";
                when x"16D9" => data <= "0110111111";
                when x"16DA" => data <= "0001100111";
                when x"16DB" => data <= "0101000100";
                when x"16DC" => data <= "1011000000";
                when x"16DD" => data <= "1111010110";
                when x"16DE" => data <= "1011110101";
                when x"16DF" => data <= "1100110111";
                when x"16E0" => data <= "0000001101";
                when x"16E1" => data <= "1010101010";
                when x"16E2" => data <= "1000010100";
                when x"16E3" => data <= "1011000000";
                when x"16E4" => data <= "0001100111";
                when x"16E5" => data <= "0110100101";
                when x"16E6" => data <= "0111111010";
                when x"16E7" => data <= "0101000100";
                when x"16E8" => data <= "1011000000";
                when x"16E9" => data <= "1000010100";
                when x"16EA" => data <= "1111010110";
                when x"16EB" => data <= "1011110101";
                when x"16EC" => data <= "0001010010";
                when x"16ED" => data <= "0010110011";
                when x"16EE" => data <= "0000001101";
                when x"16EF" => data <= "0001010010";
                when x"16F0" => data <= "1000100001";
                when x"16F1" => data <= "1111010110";
                when x"16F2" => data <= "0101000100";
                when x"16F3" => data <= "0101000100";
                when x"16F4" => data <= "0101000100";
                when x"16F5" => data <= "0001010010";
                when x"16F6" => data <= "1000100001";
                when x"16F7" => data <= "1011000000";
                when x"16F8" => data <= "0101110001";
                when x"16F9" => data <= "0001010010";
                when x"16FA" => data <= "1111010110";
                when x"16FB" => data <= "0000001101";
                when x"16FC" => data <= "1100110111";
                when x"16FD" => data <= "1011000000";
                when x"16FE" => data <= "1010101010";
                when x"16FF" => data <= "0001100111";
                when x"1700" => data <= "1010011111";
                when x"1701" => data <= "0101000100";
                when x"1702" => data <= "0001100111";
                when x"1703" => data <= "1111010110";
                when x"1704" => data <= "0001100111";
                when x"1705" => data <= "0101000100";
                when x"1706" => data <= "1100110111";
                when x"1707" => data <= "1111010110";
                when x"1708" => data <= "1111010110";
                when x"1709" => data <= "1111010110";
                when x"170A" => data <= "1011000000";
                when x"170B" => data <= "0101000100";
                when x"170C" => data <= "1011000000";
                when x"170D" => data <= "1000010100";
                when x"170E" => data <= "1010001000";
                when x"170F" => data <= "1010001000";
                when x"1710" => data <= "0001000101";
                when x"1711" => data <= "1010001000";
                when x"1712" => data <= "1010001000";
                when x"1713" => data <= "1101111111";
                when x"1714" => data <= "1101111111";
                when x"1715" => data <= "1101111111";
                when x"1716" => data <= "1101111111";
                when x"1717" => data <= "1101111111";
                when x"1718" => data <= "1110011110";
                when x"1719" => data <= "1011010111";
                when x"171A" => data <= "1010111101";
                when x"171B" => data <= "0011111011";
                when x"171C" => data <= "1101111111";
                when x"171D" => data <= "1101111111";
                when x"171E" => data <= "1101111111";
                when x"171F" => data <= "1010111101";
                when x"1720" => data <= "1101111111";
                when x"1721" => data <= "0100001100";
                when x"1722" => data <= "1101111111";
                when x"1723" => data <= "1101111111";
                when x"1724" => data <= "1000110110";
                when x"1725" => data <= "1101111111";
                when x"1726" => data <= "1011010111";
                when x"1727" => data <= "0001000101";
                when x"1728" => data <= "1101111111";
                when x"1729" => data <= "0001000101";
                when x"172A" => data <= "1101111111";
                when x"172B" => data <= "1010001000";
                when x"172C" => data <= "0110000111";
                when x"172D" => data <= "1011100010";
                when x"172E" => data <= "1100010101";
                when x"172F" => data <= "1101111111";
                when x"1730" => data <= "1101111111";
                when x"1731" => data <= "1101111111";
                when x"1732" => data <= "1101111111";
                when x"1733" => data <= "0000101111";
                when x"1734" => data <= "1101111111";
                when x"1735" => data <= "0100001100";
                when x"1736" => data <= "0011111011";
                when x"1737" => data <= "1010001000";
                when x"1738" => data <= "1101111111";
                when x"1739" => data <= "1010001000";
                when x"173A" => data <= "1101111111";
                when x"173B" => data <= "1101111111";
                when x"173C" => data <= "1101111111";
                when x"173D" => data <= "0110000111";
                when x"173E" => data <= "1101111111";
                when x"173F" => data <= "0100001100";
                when x"1740" => data <= "0001000101";
                when x"1741" => data <= "0011111011";
                when x"1742" => data <= "1101111111";
                when x"1743" => data <= "1101111111";
                when x"1744" => data <= "1101111111";
                when x"1745" => data <= "1101111111";
                when x"1746" => data <= "0111101101";
                when x"1747" => data <= "1101111111";
                when x"1748" => data <= "0111011000";
                when x"1749" => data <= "1010001000";
                when x"174A" => data <= "1011010111";
                when x"174B" => data <= "0111101101";
                when x"174C" => data <= "1010001000";
                when x"174D" => data <= "1010001000";
                when x"174E" => data <= "1100010101";
                when x"174F" => data <= "1101111111";
                when x"1750" => data <= "1010001000";
                when x"1751" => data <= "1101111111";
                when x"1752" => data <= "1010001000";
                when x"1753" => data <= "0000101111";
                when x"1754" => data <= "1101111111";
                when x"1755" => data <= "1101111111";
                when x"1756" => data <= "1101111111";
                when x"1757" => data <= "1010001000";
                when x"1758" => data <= "0011111011";
                when x"1759" => data <= "1101111111";
                when x"175A" => data <= "1010001000";
                when x"175B" => data <= "1010111101";
                when x"175C" => data <= "0000000000";
                when x"175D" => data <= "0000000000";
                when x"175E" => data <= "0000000000";
                when x"175F" => data <= "0000000000";
                when x"1760" => data <= "0000000000";
                when x"1761" => data <= "0000000000";
                when x"1762" => data <= "0000000000";
                when x"1763" => data <= "0000000000";
                when x"1764" => data <= "0000000000";
                when x"1765" => data <= "0000000000";
                when x"1766" => data <= "0000000000";
                when x"1767" => data <= "0000000000";
                when x"1768" => data <= "0000000000";
                when x"1769" => data <= "0000000000";
                when x"176A" => data <= "0000000000";
                when x"176B" => data <= "0000000000";
                when x"176C" => data <= "0000000000";
                when x"176D" => data <= "0000000000";
                when x"176E" => data <= "0000000000";
                when x"176F" => data <= "0000000000";
                when x"1770" => data <= "0000000000";
                when x"1771" => data <= "0000000000";
                when x"1772" => data <= "0000000000";
                when x"1773" => data <= "0000000000";
                when x"1774" => data <= "0000000000";
                when x"1775" => data <= "0000000000";
                when x"1776" => data <= "0000000000";
                when x"1777" => data <= "0000000000";
                when x"1778" => data <= "0000000000";
                when x"1779" => data <= "0000000000";
                when x"177A" => data <= "0000000000";
                when x"177B" => data <= "0000000000";
                when x"177C" => data <= "0000000000";
                when x"177D" => data <= "0000000000";
                when x"177E" => data <= "0000000000";
                when x"177F" => data <= "0000000000";
                when x"1780" => data <= "0000000000";
                when x"1781" => data <= "0000000000";
                when x"1782" => data <= "0000000000";
                when x"1783" => data <= "0000000000";
                when x"1784" => data <= "0000000000";
                when x"1785" => data <= "0000000000";
                when x"1786" => data <= "0000000000";
                when x"1787" => data <= "1111011011";
                when x"1788" => data <= "0000000000";
                when x"1789" => data <= "0000000000";
                when x"178A" => data <= "0000000000";
                when x"178B" => data <= "0000000000";
                when x"178C" => data <= "0000000000";
                when x"178D" => data <= "0000000000";
                when x"178E" => data <= "0000000000";
                when x"178F" => data <= "0000000000";
                when x"1790" => data <= "0000000000";
                when x"1791" => data <= "0000000000";
                when x"1792" => data <= "0000000000";
                when x"1793" => data <= "0000000000";
                when x"1794" => data <= "0000000000";
                when x"1795" => data <= "0000000000";
                when x"1796" => data <= "0000000000";
                when x"1797" => data <= "0000000000";
                when x"1798" => data <= "0000000000";
                when x"1799" => data <= "0000000000";
                when x"179A" => data <= "0000000000";
                when x"179B" => data <= "0000000000";
                when x"179C" => data <= "0000000000";
                when x"179D" => data <= "0111110111";
                when x"179E" => data <= "0000000000";
                when x"179F" => data <= "0000000000";
                when x"17A0" => data <= "0000000000";
                when x"17A1" => data <= "0000000000";
                when x"17A2" => data <= "0000000000";
                when x"17A3" => data <= "0000000000";
                when x"17A4" => data <= "0000000000";
                when x"17A5" => data <= "0000000000";
                when x"17A6" => data <= "0000000000";
                when x"17A7" => data <= "0000000000";
                when x"17A8" => data <= "0000000000";
                when x"17A9" => data <= "0000000000";
                when x"17AA" => data <= "0000000000";
                when x"17AB" => data <= "0000000000";
                when x"17AC" => data <= "0000000000";
                when x"17AD" => data <= "0000000000";
                when x"17AE" => data <= "0000000000";
                when x"17AF" => data <= "0000000000";
                when x"17B0" => data <= "0000000000";
                when x"17B1" => data <= "0000000000";
                when x"17B2" => data <= "0000000000";
                when x"17B3" => data <= "0000000000";
                when x"17B4" => data <= "0000000000";
                when x"17B5" => data <= "0000000000";
                when x"17B6" => data <= "0000000000";
                when x"17B7" => data <= "0000000000";
                when x"17B8" => data <= "0000000000";
                when x"17B9" => data <= "0000000000";
                when x"17BA" => data <= "0000000000";
                when x"17BB" => data <= "0000000000";
                when x"17BC" => data <= "0000000000";
                when x"17BD" => data <= "0000000000";
                when x"17BE" => data <= "0000000000";
                when x"17BF" => data <= "0000000000";
                when x"17C0" => data <= "0000000000";
                when x"17C1" => data <= "0000000000";
                when x"17C2" => data <= "0000000000";
                when x"17C3" => data <= "0000000000";
                when x"17C4" => data <= "0000000000";
                when x"17C5" => data <= "0000000000";
                when x"17C6" => data <= "0000000000";
                when x"17C7" => data <= "0000000000";
                when x"17C8" => data <= "0000000000";
                when x"17C9" => data <= "0000000000";
                when x"17CA" => data <= "0000000000";
                when x"17CB" => data <= "0000000000";
                when x"17CC" => data <= "0000000000";
                when x"17CD" => data <= "0000000000";
                when x"17CE" => data <= "0000000000";
                when x"17CF" => data <= "0000000000";
                when x"17D0" => data <= "0000000000";
                when x"17D1" => data <= "0000000000";
                when x"17D2" => data <= "0000000000";
                when x"17D3" => data <= "0000000000";
                when x"17D4" => data <= "0000000000";
                when x"17D5" => data <= "0000000000";
                when x"17D6" => data <= "0000000000";
                when x"17D7" => data <= "0000000000";
                when x"17D8" => data <= "0000000000";
                when x"17D9" => data <= "0000000000";
                when x"17DA" => data <= "0000000000";
                when x"17DB" => data <= "0000000000";
                when x"17DC" => data <= "0000000000";
                when x"17DD" => data <= "0000000000";
                when x"17DE" => data <= "0000000000";
                when x"17DF" => data <= "0000000000";
                when x"17E0" => data <= "1011001101";
                when x"17E1" => data <= "0000000000";
                when x"17E2" => data <= "0000000000";
                when x"17E3" => data <= "0000000000";
                when x"17E4" => data <= "0000000000";
                when x"17E5" => data <= "0000000000";
                when x"17E6" => data <= "0000000000";
                when x"17E7" => data <= "0000000000";
                when x"17E8" => data <= "0000000000";
                when x"17E9" => data <= "0000000000";
                when x"17EA" => data <= "0000000000";
                when x"17EB" => data <= "0000000000";
                when x"17EC" => data <= "0000000000";
                when x"17ED" => data <= "0000000000";
                when x"17EE" => data <= "0000000000";
                when x"17EF" => data <= "0000000000";
                when x"17F0" => data <= "0000000000";
                when x"17F1" => data <= "0000000000";
                when x"17F2" => data <= "0000000000";
                when x"17F3" => data <= "0000000000";
                when x"17F4" => data <= "0000000000";
                when x"17F5" => data <= "0000000000";
                when x"17F6" => data <= "0000000000";
                when x"17F7" => data <= "0000000000";
                when x"17F8" => data <= "0000000000";
                when x"17F9" => data <= "0000000000";
                when x"17FA" => data <= "0000000000";
                when x"17FB" => data <= "0000000000";
                when x"17FC" => data <= "0000000000";
                when x"17FD" => data <= "0000000000";
                when x"17FE" => data <= "0000000000";
                when x"17FF" => data <= "0000000000";
                when x"1800" => data <= "0000000000";
                when x"1801" => data <= "0000000000";
                when x"1802" => data <= "0000000000";
                when x"1803" => data <= "0000000000";
                when x"1804" => data <= "0000000000";
                when x"1805" => data <= "0000000000";
                when x"1806" => data <= "0000000000";
                when x"1807" => data <= "0000000000";
                when x"1808" => data <= "0000000000";
                when x"1809" => data <= "0000000000";
                when x"180A" => data <= "0000000000";
                when x"180B" => data <= "0000000000";
                when x"180C" => data <= "0000000000";
                when x"180D" => data <= "0000000000";
                when x"180E" => data <= "0000000000";
                when x"180F" => data <= "0000000000";
                when x"1810" => data <= "0000000000";
                when x"1811" => data <= "0000000000";
                when x"1812" => data <= "0000000000";
                when x"1813" => data <= "0000000000";
                when x"1814" => data <= "0000000000";
                when x"1815" => data <= "0000000000";
                when x"1816" => data <= "0000000000";
                when x"1817" => data <= "0000000000";
                when x"1818" => data <= "0000000000";
                when x"1819" => data <= "0000000000";
                when x"181A" => data <= "0000000000";
                when x"181B" => data <= "0000000000";
                when x"181C" => data <= "0000000000";
                when x"181D" => data <= "0000000000";
                when x"181E" => data <= "0000000000";
                when x"181F" => data <= "0000000000";
                when x"1820" => data <= "0000000000";
                when x"1821" => data <= "0000000000";
                when x"1822" => data <= "0000000000";
                when x"1823" => data <= "0000000000";
                when x"1824" => data <= "0000000000";
                when x"1825" => data <= "0000000000";
                when x"1826" => data <= "0000000000";
                when x"1827" => data <= "0000000000";
                when x"1828" => data <= "0000000000";
                when x"1829" => data <= "0000000000";
                when x"182A" => data <= "0000000000";
                when x"182B" => data <= "0000000000";
                when x"182C" => data <= "0000000000";
                when x"182D" => data <= "0000000000";
                when x"182E" => data <= "0000000000";
                when x"182F" => data <= "0000000000";
                when x"1830" => data <= "0000000000";
                when x"1831" => data <= "0000000000";
                when x"1832" => data <= "0000000000";
                when x"1833" => data <= "0000000000";
                when x"1834" => data <= "0000000000";
                when x"1835" => data <= "0000000000";
                when x"1836" => data <= "0000000000";
                when x"1837" => data <= "0000000000";
                when x"1838" => data <= "0100010110";
                when x"1839" => data <= "0000000000";
                when x"183A" => data <= "0000000000";
                when x"183B" => data <= "0000000000";
                when x"183C" => data <= "0000000000";
                when x"183D" => data <= "0000000000";
                when x"183E" => data <= "0000000000";
                when x"183F" => data <= "0000000000";
                when x"1840" => data <= "0000000000";
                when x"1841" => data <= "0000000000";
                when x"1842" => data <= "0000000000";
                when x"1843" => data <= "0000000000";
                when x"1844" => data <= "0000000000";
                when x"1845" => data <= "0000000000";
                when x"1846" => data <= "0000000000";
                when x"1847" => data <= "0000000000";
                when x"1848" => data <= "0000000000";
                when x"1849" => data <= "0000000000";
                when x"184A" => data <= "0000000000";
                when x"184B" => data <= "0000000000";
                when x"184C" => data <= "0000000000";
                when x"184D" => data <= "0000000000";
                when x"184E" => data <= "0000000000";
                when x"184F" => data <= "0000000000";
                when x"1850" => data <= "0000000000";
                when x"1851" => data <= "0000000000";
                when x"1852" => data <= "0000000000";
                when x"1853" => data <= "0000000000";
                when x"1854" => data <= "0000000000";
                when x"1855" => data <= "0000000000";
                when x"1856" => data <= "0000000000";
                when x"1857" => data <= "0000000000";
                when x"1858" => data <= "0000000000";
                when x"1859" => data <= "0000000000";
                when x"185A" => data <= "0000000000";
                when x"185B" => data <= "0000000000";
                when x"185C" => data <= "0000000000";
                when x"185D" => data <= "0000000000";
                when x"185E" => data <= "0000000000";
                when x"185F" => data <= "0000000000";
                when x"1860" => data <= "0000000000";
                when x"1861" => data <= "0000000000";
                when x"1862" => data <= "0000000000";
                when x"1863" => data <= "0000000000";
                when x"1864" => data <= "0000000000";
                when x"1865" => data <= "0000000000";
                when x"1866" => data <= "0000000000";
                when x"1867" => data <= "0000000000";
                when x"1868" => data <= "0000000000";
                when x"1869" => data <= "0000000000";
                when x"186A" => data <= "0000000000";
                when x"186B" => data <= "0000000000";
                when x"186C" => data <= "0000000000";
                when x"186D" => data <= "0000000000";
                when x"186E" => data <= "0000000000";
                when x"186F" => data <= "0000000000";
                when x"1870" => data <= "0000000000";
                when x"1871" => data <= "0000000000";
                when x"1872" => data <= "0000000000";
                when x"1873" => data <= "0000000000";
                when x"1874" => data <= "0000000000";
                when x"1875" => data <= "0000000000";
                when x"1876" => data <= "0000000000";
                when x"1877" => data <= "0000000000";
                when x"1878" => data <= "0000000000";
                when x"1879" => data <= "0000000000";
                when x"187A" => data <= "0000000000";
                when x"187B" => data <= "0000000000";
                when x"187C" => data <= "0000000000";
                when x"187D" => data <= "0000000000";
                when x"187E" => data <= "0000000000";
                when x"187F" => data <= "0000000000";
                when x"1880" => data <= "0000000000";
                when x"1881" => data <= "0000000000";
                when x"1882" => data <= "0000000000";
                when x"1883" => data <= "0000000000";
                when x"1884" => data <= "0000000000";
                when x"1885" => data <= "0000000000";
                when x"1886" => data <= "0000000000";
                when x"1887" => data <= "0000000000";
                when x"1888" => data <= "0000000000";
                when x"1889" => data <= "0000000000";
                when x"188A" => data <= "0000000000";
                when x"188B" => data <= "0000000000";
                when x"188C" => data <= "0000000000";
                when x"188D" => data <= "0000000000";
                when x"188E" => data <= "0000000000";
                when x"188F" => data <= "0000000000";
                when x"1890" => data <= "0000000000";
                when x"1891" => data <= "0000000000";
                when x"1892" => data <= "0000000000";
                when x"1893" => data <= "0000000000";
                when x"1894" => data <= "0000000000";
                when x"1895" => data <= "0000000000";
                when x"1896" => data <= "0000000000";
                when x"1897" => data <= "0000000000";
                when x"1898" => data <= "0000000000";
                when x"1899" => data <= "0000000000";
                when x"189A" => data <= "0000000000";
                when x"189B" => data <= "0000000000";
                when x"189C" => data <= "0000000000";
                when x"189D" => data <= "0000000000";
                when x"189E" => data <= "0000000000";
                when x"189F" => data <= "0000000000";
                when x"18A0" => data <= "0000000000";
                when x"18A1" => data <= "0000000000";
                when x"18A2" => data <= "0000000000";
                when x"18A3" => data <= "0000000000";
                when x"18A4" => data <= "0000000000";
                when x"18A5" => data <= "0000000000";
                when x"18A6" => data <= "0000000000";
                when x"18A7" => data <= "0000000000";
                when x"18A8" => data <= "0000000000";
                when x"18A9" => data <= "0000000000";
                when x"18AA" => data <= "0000000000";
                when x"18AB" => data <= "0000000000";
                when x"18AC" => data <= "0000000000";
                when x"18AD" => data <= "0000000000";
                when x"18AE" => data <= "0000000000";
                when x"18AF" => data <= "0000000000";
                when x"18B0" => data <= "0000000000";
                when x"18B1" => data <= "0000000000";
                when x"18B2" => data <= "0000000000";
                when x"18B3" => data <= "0000000000";
                when x"18B4" => data <= "0000000000";
                when x"18B5" => data <= "0000000000";
                when x"18B6" => data <= "0000000000";
                when x"18B7" => data <= "0000000000";
                when x"18B8" => data <= "0000000000";
                when x"18B9" => data <= "0000000000";
                when x"18BA" => data <= "0000000000";
                when x"18BB" => data <= "0000000000";
                when x"18BC" => data <= "0000000000";
                when x"18BD" => data <= "0000000000";
                when x"18BE" => data <= "0000000000";
                when x"18BF" => data <= "0000000000";
                when x"18C0" => data <= "0000000000";
                when x"18C1" => data <= "0000000000";
                when x"18C2" => data <= "0000000000";
                when x"18C3" => data <= "0000000000";
                when x"18C4" => data <= "0000000000";
                when x"18C5" => data <= "0000000000";
                when x"18C6" => data <= "0000000000";
                when x"18C7" => data <= "0000000000";
                when x"18C8" => data <= "0000000000";
                when x"18C9" => data <= "0000000000";
                when x"18CA" => data <= "0000000000";
                when x"18CB" => data <= "0000000000";
                when x"18CC" => data <= "0000000000";
                when x"18CD" => data <= "0000000000";
                when x"18CE" => data <= "0000000000";
                when x"18CF" => data <= "0000000000";
                when x"18D0" => data <= "0000000000";
                when x"18D1" => data <= "0000000000";
                when x"18D2" => data <= "0000000000";
                when x"18D3" => data <= "0000000000";
                when x"18D4" => data <= "0000000000";
                when x"18D5" => data <= "0000000000";
                when x"18D6" => data <= "0000000000";
                when x"18D7" => data <= "0000000000";
                when x"18D8" => data <= "0000000000";
                when x"18D9" => data <= "0000000000";
                when x"18DA" => data <= "0000000000";
                when x"18DB" => data <= "0000000000";
                when x"18DC" => data <= "0000000000";
                when x"18DD" => data <= "0000000000";
                when x"18DE" => data <= "0000000000";
                when x"18DF" => data <= "0000000000";
                when x"18E0" => data <= "0000000000";
                when x"18E1" => data <= "0000000000";
                when x"18E2" => data <= "0000000000";
                when x"18E3" => data <= "0000000000";
                when x"18E4" => data <= "0000000000";
                when x"18E5" => data <= "0000000000";
                when x"18E6" => data <= "0000000000";
                when x"18E7" => data <= "0000000000";
                when x"18E8" => data <= "0000000000";
                when x"18E9" => data <= "0000000000";
                when x"18EA" => data <= "0000000000";
                when x"18EB" => data <= "0000000000";
                when x"18EC" => data <= "0000000000";
                when x"18ED" => data <= "0000000000";
                when x"18EE" => data <= "0000000000";
                when x"18EF" => data <= "0000000000";
                when x"18F0" => data <= "0000000000";
                when x"18F1" => data <= "0000000000";
                when x"18F2" => data <= "0000000000";
                when x"18F3" => data <= "0000000000";
                when x"18F4" => data <= "0000000000";
                when x"18F5" => data <= "0000000000";
                when x"18F6" => data <= "0000000000";
                when x"18F7" => data <= "0000000000";
                when x"18F8" => data <= "0000000000";
                when x"18F9" => data <= "0000000000";
                when x"18FA" => data <= "0000000000";
                when x"18FB" => data <= "0000000000";
                when x"18FC" => data <= "0000000000";
                when x"18FD" => data <= "0000000000";
                when x"18FE" => data <= "0000000000";
                when x"18FF" => data <= "0000000000";
                when x"1900" => data <= "0000000000";
                when x"1901" => data <= "0000000000";
                when x"1902" => data <= "0000000000";
                when x"1903" => data <= "0000000000";
                when x"1904" => data <= "0000000000";
                when x"1905" => data <= "0000000000";
                when x"1906" => data <= "0000000000";
                when x"1907" => data <= "0000000000";
                when x"1908" => data <= "0000000000";
                when x"1909" => data <= "0000000000";
                when x"190A" => data <= "0000000000";
                when x"190B" => data <= "0000000000";
                when x"190C" => data <= "0000000000";
                when x"190D" => data <= "0000000000";
                when x"190E" => data <= "0000000000";
                when x"190F" => data <= "0000000000";
                when x"1910" => data <= "0000000000";
                when x"1911" => data <= "0000000000";
                when x"1912" => data <= "0000000000";
                when x"1913" => data <= "0000000000";
                when x"1914" => data <= "0000000000";
                when x"1915" => data <= "0000000000";
                when x"1916" => data <= "0000000000";
                when x"1917" => data <= "0000000000";
                when x"1918" => data <= "0000000000";
                when x"1919" => data <= "0000000000";
                when x"191A" => data <= "0000000000";
                when x"191B" => data <= "0000000000";
                when x"191C" => data <= "0000000000";
                when x"191D" => data <= "0000000000";
                when x"191E" => data <= "0000000000";
                when x"191F" => data <= "0000000000";
                when x"1920" => data <= "0000000000";
                when x"1921" => data <= "0000000000";
                when x"1922" => data <= "0000000000";
                when x"1923" => data <= "0000000000";
                when x"1924" => data <= "0000000000";
                when x"1925" => data <= "0000000000";
                when x"1926" => data <= "0111110111";
                when x"1927" => data <= "0000000000";
                when x"1928" => data <= "0000000000";
                when x"1929" => data <= "0000000000";
                when x"192A" => data <= "0000000000";
                when x"192B" => data <= "0000000000";
                when x"192C" => data <= "0000000000";
                when x"192D" => data <= "0000000000";
                when x"192E" => data <= "0000000000";
                when x"192F" => data <= "0000000000";
                when x"1930" => data <= "0000000000";
                when x"1931" => data <= "0000000000";
                when x"1932" => data <= "0000000000";
                when x"1933" => data <= "0000000000";
                when x"1934" => data <= "0000000000";
                when x"1935" => data <= "0000000000";
                when x"1936" => data <= "0000000000";
                when x"1937" => data <= "0000000000";
                when x"1938" => data <= "0000000000";
                when x"1939" => data <= "0000000000";
                when x"193A" => data <= "0000000000";
                when x"193B" => data <= "0000000000";
                when x"193C" => data <= "0000000000";
                when x"193D" => data <= "0000000000";
                when x"193E" => data <= "0000000000";
                when x"193F" => data <= "0000000000";
                when x"1940" => data <= "0000000000";
                when x"1941" => data <= "0000000000";
                when x"1942" => data <= "0000000000";
                when x"1943" => data <= "0000000000";
                when x"1944" => data <= "0000000000";
                when x"1945" => data <= "0000000000";
                when x"1946" => data <= "0000000000";
                when x"1947" => data <= "0000000000";
                when x"1948" => data <= "0000000000";
                when x"1949" => data <= "0000000000";
                when x"194A" => data <= "0000000000";
                when x"194B" => data <= "0000000000";
                when x"194C" => data <= "0000000000";
                when x"194D" => data <= "0000000000";
                when x"194E" => data <= "0000000000";
                when x"194F" => data <= "0000000000";
                when x"1950" => data <= "0000000000";
                when x"1951" => data <= "0000000000";
                when x"1952" => data <= "0000000000";
                when x"1953" => data <= "0000000000";
                when x"1954" => data <= "0000000000";
                when x"1955" => data <= "0000000000";
                when x"1956" => data <= "0000000000";
                when x"1957" => data <= "0000000000";
                when x"1958" => data <= "0000000000";
                when x"1959" => data <= "0000000000";
                when x"195A" => data <= "0000000000";
                when x"195B" => data <= "0000000000";
                when x"195C" => data <= "0000000000";
                when x"195D" => data <= "0000000000";
                when x"195E" => data <= "0000000000";
                when x"195F" => data <= "0000000000";
                when x"1960" => data <= "0000000000";
                when x"1961" => data <= "0000000000";
                when x"1962" => data <= "0000000000";
                when x"1963" => data <= "0000000000";
                when x"1964" => data <= "0000000000";
                when x"1965" => data <= "0000000000";
                when x"1966" => data <= "0000000000";
                when x"1967" => data <= "0000000000";
                when x"1968" => data <= "0000000000";
                when x"1969" => data <= "0000000000";
                when x"196A" => data <= "0000000000";
                when x"196B" => data <= "0000000000";
                when x"196C" => data <= "0000000000";
                when x"196D" => data <= "0000000000";
                when x"196E" => data <= "0000000000";
                when x"196F" => data <= "0000000000";
                when x"1970" => data <= "0000000000";
                when x"1971" => data <= "0000000000";
                when x"1972" => data <= "0000000000";
                when x"1973" => data <= "0000000000";
                when x"1974" => data <= "0000000000";
                when x"1975" => data <= "0000000000";
                when x"1976" => data <= "0000000000";
                when x"1977" => data <= "0000000000";
                when x"1978" => data <= "0000000000";
                when x"1979" => data <= "0000000000";
                when x"197A" => data <= "0000000000";
                when x"197B" => data <= "0000000000";
                when x"197C" => data <= "0000000000";
                when x"197D" => data <= "0000000000";
                when x"197E" => data <= "0000000000";
                when x"197F" => data <= "0000000000";
                when x"1980" => data <= "0000000000";
                when x"1981" => data <= "0000000000";
                when x"1982" => data <= "0000000000";
                when x"1983" => data <= "0000000000";
                when x"1984" => data <= "0000000000";
                when x"1985" => data <= "0000000000";
                when x"1986" => data <= "0000000000";
                when x"1987" => data <= "0000000000";
                when x"1988" => data <= "0000000000";
                when x"1989" => data <= "0000000000";
                when x"198A" => data <= "0000000000";
                when x"198B" => data <= "0000000000";
                when x"198C" => data <= "0000000000";
                when x"198D" => data <= "0000000000";
                when x"198E" => data <= "0000000000";
                when x"198F" => data <= "0000000000";
                when x"1990" => data <= "0000000000";
                when x"1991" => data <= "0000000000";
                when x"1992" => data <= "0000000000";
                when x"1993" => data <= "0000000000";
                when x"1994" => data <= "0000000000";
                when x"1995" => data <= "0000000000";
                when x"1996" => data <= "0000000000";
                when x"1997" => data <= "0000000000";
                when x"1998" => data <= "0000000000";
                when x"1999" => data <= "0000000000";
                when x"199A" => data <= "0000000000";
                when x"199B" => data <= "0000000000";
                when x"199C" => data <= "0000000000";
                when x"199D" => data <= "0000000000";
                when x"199E" => data <= "0000000000";
                when x"199F" => data <= "0000000000";
                when x"19A0" => data <= "0000000000";
                when x"19A1" => data <= "0000000000";
                when x"19A2" => data <= "0000000000";
                when x"19A3" => data <= "0000000000";
                when x"19A4" => data <= "0000000000";
                when x"19A5" => data <= "0000000000";
                when x"19A6" => data <= "0000000000";
                when x"19A7" => data <= "0000000000";
                when x"19A8" => data <= "0000000000";
                when x"19A9" => data <= "0000000000";
                when x"19AA" => data <= "0000000000";
                when x"19AB" => data <= "0000000000";
                when x"19AC" => data <= "0000000000";
                when x"19AD" => data <= "0000000000";
                when x"19AE" => data <= "0000000000";
                when x"19AF" => data <= "0000000000";
                when x"19B0" => data <= "0000000000";
                when x"19B1" => data <= "0000000000";
                when x"19B2" => data <= "0000000000";
                when x"19B3" => data <= "0000000000";
                when x"19B4" => data <= "0000000000";
                when x"19B5" => data <= "0000000000";
                when x"19B6" => data <= "0000000000";
                when x"19B7" => data <= "0000000000";
                when x"19B8" => data <= "0000000000";
                when x"19B9" => data <= "0000000000";
                when x"19BA" => data <= "0000000000";
                when x"19BB" => data <= "0000000000";
                when x"19BC" => data <= "0000000000";
                when x"19BD" => data <= "0000000000";
                when x"19BE" => data <= "0000000000";
                when x"19BF" => data <= "0000000000";
                when x"19C0" => data <= "0000000000";
                when x"19C1" => data <= "0000000000";
                when x"19C2" => data <= "0000000000";
                when x"19C3" => data <= "0000000000";
                when x"19C4" => data <= "0000000000";
                when x"19C5" => data <= "0000000000";
                when x"19C6" => data <= "0000000000";
                when x"19C7" => data <= "0000000000";
                when x"19C8" => data <= "0000000000";
                when x"19C9" => data <= "0000000000";
                when x"19CA" => data <= "0000000000";
                when x"19CB" => data <= "0000000000";
                when x"19CC" => data <= "0000000000";
                when x"19CD" => data <= "0000000000";
                when x"19CE" => data <= "0000000000";
                when x"19CF" => data <= "0000000000";
                when x"19D0" => data <= "0000000000";
                when x"19D1" => data <= "0000000000";
                when x"19D2" => data <= "0000000000";
                when x"19D3" => data <= "0000000000";
                when x"19D4" => data <= "0000000000";
                when x"19D5" => data <= "0000000000";
                when x"19D6" => data <= "0000000000";
                when x"19D7" => data <= "0000000000";
                when x"19D8" => data <= "0000000000";
                when x"19D9" => data <= "0000000000";
                when x"19DA" => data <= "0000000000";
                when x"19DB" => data <= "0000000000";
                when x"19DC" => data <= "0000000000";
                when x"19DD" => data <= "0000000000";
                when x"19DE" => data <= "0000000000";
                when x"19DF" => data <= "0000000000";
                when x"19E0" => data <= "0000000000";
                when x"19E1" => data <= "0000000000";
                when x"19E2" => data <= "0000000000";
                when x"19E3" => data <= "0000000000";
                when x"19E4" => data <= "0000000000";
                when x"19E5" => data <= "0000000000";
                when x"19E6" => data <= "0000000000";
                when x"19E7" => data <= "0000000000";
                when x"19E8" => data <= "0000000000";
                when x"19E9" => data <= "0000000000";
                when x"19EA" => data <= "0000000000";
                when x"19EB" => data <= "0000000000";
                when x"19EC" => data <= "0000000000";
                when x"19ED" => data <= "0000000000";
                when x"19EE" => data <= "0000000000";
                when x"19EF" => data <= "0000000000";
                when x"19F0" => data <= "0000000000";
                when x"19F1" => data <= "0000000000";
                when x"19F2" => data <= "0000000000";
                when x"19F3" => data <= "0000000000";
                when x"19F4" => data <= "0000000000";
                when x"19F5" => data <= "0000000000";
                when x"19F6" => data <= "0000000000";
                when x"19F7" => data <= "0000000000";
                when x"19F8" => data <= "0000000000";
                when x"19F9" => data <= "0000000000";
                when x"19FA" => data <= "0000000000";
                when x"19FB" => data <= "0000000000";
                when x"19FC" => data <= "0000000000";
                when x"19FD" => data <= "0000000000";
                when x"19FE" => data <= "0000000000";
                when x"19FF" => data <= "0000000000";
                when x"1A00" => data <= "0000000000";
                when x"1A01" => data <= "0000000000";
                when x"1A02" => data <= "0000000000";
                when x"1A03" => data <= "0000000000";
                when x"1A04" => data <= "0000000000";
                when x"1A05" => data <= "0000000000";
                when x"1A06" => data <= "0000000000";
                when x"1A07" => data <= "0000000000";
                when x"1A08" => data <= "0000000000";
                when x"1A09" => data <= "0000000000";
                when x"1A0A" => data <= "0000000000";
                when x"1A0B" => data <= "0000000000";
                when x"1A0C" => data <= "0000000000";
                when x"1A0D" => data <= "0000000000";
                when x"1A0E" => data <= "0000000000";
                when x"1A0F" => data <= "0000000000";
                when x"1A10" => data <= "0000000000";
                when x"1A11" => data <= "0000000000";
                when x"1A12" => data <= "0000000000";
                when x"1A13" => data <= "0000000000";
                when x"1A14" => data <= "0000000000";
                when x"1A15" => data <= "0000000000";
                when x"1A16" => data <= "0000000000";
                when x"1A17" => data <= "0000000000";
                when x"1A18" => data <= "0000000000";
                when x"1A19" => data <= "0000000000";
                when x"1A1A" => data <= "0000000000";
                when x"1A1B" => data <= "0000000000";
                when x"1A1C" => data <= "0000000000";
                when x"1A1D" => data <= "0000000000";
                when x"1A1E" => data <= "0000000000";
                when x"1A1F" => data <= "0000000000";
                when x"1A20" => data <= "0000000000";
                when x"1A21" => data <= "0000000000";
                when x"1A22" => data <= "0000000000";
                when x"1A23" => data <= "0000000000";
                when x"1A24" => data <= "0000000000";
                when x"1A25" => data <= "0000000000";
                when x"1A26" => data <= "0000000000";
                when x"1A27" => data <= "0000000000";
                when x"1A28" => data <= "0000000000";
                when x"1A29" => data <= "0000000000";
                when x"1A2A" => data <= "0000000000";
                when x"1A2B" => data <= "0000000000";
                when x"1A2C" => data <= "0000000000";
                when x"1A2D" => data <= "0000000000";
                when x"1A2E" => data <= "0000000000";
                when x"1A2F" => data <= "0000000000";
                when x"1A30" => data <= "0000000000";
                when x"1A31" => data <= "0000000000";
                when x"1A32" => data <= "0000000000";
                when x"1A33" => data <= "0000000000";
                when x"1A34" => data <= "0000000000";
                when x"1A35" => data <= "0000000000";
                when x"1A36" => data <= "0000000000";
                when x"1A37" => data <= "0000000000";
                when x"1A38" => data <= "0000000000";
                when x"1A39" => data <= "0000000000";
                when x"1A3A" => data <= "0000000000";
                when x"1A3B" => data <= "0000000000";
                when x"1A3C" => data <= "0000000000";
                when x"1A3D" => data <= "0000000000";
                when x"1A3E" => data <= "0000000000";
                when x"1A3F" => data <= "0000000000";
                when x"1A40" => data <= "0000000000";
                when x"1A41" => data <= "0000000000";
                when x"1A42" => data <= "0000000000";
                when x"1A43" => data <= "0000000000";
                when x"1A44" => data <= "0000000000";
                when x"1A45" => data <= "0000000000";
                when x"1A46" => data <= "0000000000";
                when x"1A47" => data <= "0000000000";
                when x"1A48" => data <= "0000000000";
                when x"1A49" => data <= "0000000000";
                when x"1A4A" => data <= "0000000000";
                when x"1A4B" => data <= "0000000000";
                when x"1A4C" => data <= "0000000000";
                when x"1A4D" => data <= "0000000000";
                when x"1A4E" => data <= "0000000000";
                when x"1A4F" => data <= "0000000000";
                when x"1A50" => data <= "0000000000";
                when x"1A51" => data <= "0000000000";
                when x"1A52" => data <= "0000000000";
                when x"1A53" => data <= "0000000000";
                when x"1A54" => data <= "0000000000";
                when x"1A55" => data <= "0000000000";
                when x"1A56" => data <= "0000000000";
                when x"1A57" => data <= "0000000000";
                when x"1A58" => data <= "0000000000";
                when x"1A59" => data <= "0000000000";
                when x"1A5A" => data <= "0000000000";
                when x"1A5B" => data <= "0000000000";
                when x"1A5C" => data <= "0000000000";
                when x"1A5D" => data <= "0000000000";
                when x"1A5E" => data <= "0000000000";
                when x"1A5F" => data <= "0000000000";
                when x"1A60" => data <= "0000000000";
                when x"1A61" => data <= "0000000000";
                when x"1A62" => data <= "0000000000";
                when x"1A63" => data <= "0000000000";
                when x"1A64" => data <= "0000000000";
                when x"1A65" => data <= "0000000000";
                when x"1A66" => data <= "0000000000";
                when x"1A67" => data <= "0000000000";
                when x"1A68" => data <= "0000000000";
                when x"1A69" => data <= "0000000000";
                when x"1A6A" => data <= "0000000000";
                when x"1A6B" => data <= "0000000000";
                when x"1A6C" => data <= "0000000000";
                when x"1A6D" => data <= "0000000000";
                when x"1A6E" => data <= "0000000000";
                when x"1A6F" => data <= "0000000000";
                when x"1A70" => data <= "0000000000";
                when x"1A71" => data <= "0000000000";
                when x"1A72" => data <= "0000000000";
                when x"1A73" => data <= "0000000000";
                when x"1A74" => data <= "0000000000";
                when x"1A75" => data <= "0000000000";
                when x"1A76" => data <= "0000000000";
                when x"1A77" => data <= "0000000000";
                when x"1A78" => data <= "0000000000";
                when x"1A79" => data <= "0000000000";
                when x"1A7A" => data <= "0000000000";
                when x"1A7B" => data <= "0000000000";
                when x"1A7C" => data <= "0000000000";
                when x"1A7D" => data <= "0000000000";
                when x"1A7E" => data <= "0000000000";
                when x"1A7F" => data <= "0000000000";
                when x"1A80" => data <= "0000000000";
                when x"1A81" => data <= "0000000000";
                when x"1A82" => data <= "0000000000";
                when x"1A83" => data <= "0000000000";
                when x"1A84" => data <= "0000000000";
                when x"1A85" => data <= "0000000000";
                when x"1A86" => data <= "0000000000";
                when x"1A87" => data <= "0000000000";
                when x"1A88" => data <= "0000000000";
                when x"1A89" => data <= "0000000000";
                when x"1A8A" => data <= "0000000000";
                when x"1A8B" => data <= "0000000000";
                when x"1A8C" => data <= "0000000000";
                when x"1A8D" => data <= "0000000000";
                when x"1A8E" => data <= "0000000000";
                when x"1A8F" => data <= "0000000000";
                when x"1A90" => data <= "0000000000";
                when x"1A91" => data <= "0000000000";
                when x"1A92" => data <= "0000000000";
                when x"1A93" => data <= "0000000000";
                when x"1A94" => data <= "0000000000";
                when x"1A95" => data <= "0000000000";
                when x"1A96" => data <= "0000000000";
                when x"1A97" => data <= "0000000000";
                when x"1A98" => data <= "0000000000";
                when x"1A99" => data <= "0000000000";
                when x"1A9A" => data <= "0000000000";
                when x"1A9B" => data <= "0000000000";
                when x"1A9C" => data <= "0000000000";
                when x"1A9D" => data <= "0000000000";
                when x"1A9E" => data <= "0000000000";
                when x"1A9F" => data <= "0000000000";
                when x"1AA0" => data <= "0000000000";
                when x"1AA1" => data <= "0000000000";
                when x"1AA2" => data <= "0000000000";
                when x"1AA3" => data <= "0000000000";
                when x"1AA4" => data <= "0000000000";
                when x"1AA5" => data <= "0000000000";
                when x"1AA6" => data <= "0000000000";
                when x"1AA7" => data <= "0000000000";
                when x"1AA8" => data <= "0000000000";
                when x"1AA9" => data <= "0000000000";
                when x"1AAA" => data <= "0000000000";
                when x"1AAB" => data <= "0000000000";
                when x"1AAC" => data <= "0000000000";
                when x"1AAD" => data <= "0000000000";
                when x"1AAE" => data <= "0000000000";
                when x"1AAF" => data <= "0000000000";
                when x"1AB0" => data <= "0000000000";
                when x"1AB1" => data <= "0000000000";
                when x"1AB2" => data <= "0000000000";
                when x"1AB3" => data <= "0000000000";
                when x"1AB4" => data <= "0000000000";
                when x"1AB5" => data <= "0000000000";
                when x"1AB6" => data <= "0000000000";
                when x"1AB7" => data <= "0000000000";
                when x"1AB8" => data <= "0000000000";
                when x"1AB9" => data <= "0000000000";
                when x"1ABA" => data <= "0000000000";
                when x"1ABB" => data <= "0000000000";
                when x"1ABC" => data <= "0000000000";
                when x"1ABD" => data <= "0000000000";
                when x"1ABE" => data <= "0000000000";
                when x"1ABF" => data <= "0000000000";
                when x"1AC0" => data <= "0000000000";
                when x"1AC1" => data <= "0000000000";
                when x"1AC2" => data <= "0000000000";
                when x"1AC3" => data <= "0000000000";
                when x"1AC4" => data <= "0000000000";
                when x"1AC5" => data <= "0000000000";
                when x"1AC6" => data <= "0000000000";
                when x"1AC7" => data <= "0000000000";
                when x"1AC8" => data <= "0000000000";
                when x"1AC9" => data <= "0000000000";
                when x"1ACA" => data <= "0000000000";
                when x"1ACB" => data <= "0000000000";
                when x"1ACC" => data <= "0000000000";
                when x"1ACD" => data <= "0000000000";
                when x"1ACE" => data <= "0000000000";
                when x"1ACF" => data <= "0000000000";
                when x"1AD0" => data <= "0000000000";
                when x"1AD1" => data <= "0000000000";
                when x"1AD2" => data <= "0000000000";
                when x"1AD3" => data <= "0000000000";
                when x"1AD4" => data <= "0000000000";
                when x"1AD5" => data <= "0000000000";
                when x"1AD6" => data <= "0000000000";
                when x"1AD7" => data <= "0000000000";
                when x"1AD8" => data <= "0000000000";
                when x"1AD9" => data <= "0000000000";
                when x"1ADA" => data <= "0000000000";
                when x"1ADB" => data <= "0000000000";
                when x"1ADC" => data <= "0000000000";
                when x"1ADD" => data <= "0000000000";
                when x"1ADE" => data <= "0000000000";
                when x"1ADF" => data <= "0000000000";
                when x"1AE0" => data <= "0000000000";
                when x"1AE1" => data <= "0000000000";
                when x"1AE2" => data <= "0000000000";
                when x"1AE3" => data <= "0000000000";
                when x"1AE4" => data <= "0000000000";
                when x"1AE5" => data <= "0000000000";
                when x"1AE6" => data <= "0000000000";
                when x"1AE7" => data <= "0000000000";
                when x"1AE8" => data <= "0000000000";
                when x"1AE9" => data <= "0000000000";
                when x"1AEA" => data <= "0000000000";
                when x"1AEB" => data <= "0000000000";
                when x"1AEC" => data <= "0000000000";
                when x"1AED" => data <= "0000000000";
                when x"1AEE" => data <= "0111110111";
                when x"1AEF" => data <= "0000000000";
                when x"1AF0" => data <= "0000000000";
                when x"1AF1" => data <= "0000000000";
                when x"1AF2" => data <= "0000000000";
                when x"1AF3" => data <= "0000000000";
                when x"1AF4" => data <= "0000000000";
                when x"1AF5" => data <= "0000000000";
                when x"1AF6" => data <= "0000000000";
                when x"1AF7" => data <= "0000000000";
                when x"1AF8" => data <= "0000000000";
                when x"1AF9" => data <= "0000000000";
                when x"1AFA" => data <= "0000000000";
                when x"1AFB" => data <= "0000000000";
                when x"1AFC" => data <= "0000000000";
                when x"1AFD" => data <= "0000000000";
                when x"1AFE" => data <= "0000000000";
                when x"1AFF" => data <= "0000000000";
                when x"1B00" => data <= "0000000000";
                when x"1B01" => data <= "0000000000";
                when x"1B02" => data <= "0000000000";
                when x"1B03" => data <= "0000000000";
                when x"1B04" => data <= "0000000000";
                when x"1B05" => data <= "0000000000";
                when x"1B06" => data <= "0000000000";
                when x"1B07" => data <= "0000000000";
                when x"1B08" => data <= "0000000000";
                when x"1B09" => data <= "0000000000";
                when x"1B0A" => data <= "0000000000";
                when x"1B0B" => data <= "0000000000";
                when x"1B0C" => data <= "0000000000";
                when x"1B0D" => data <= "0000000000";
                when x"1B0E" => data <= "0000000000";
                when x"1B0F" => data <= "0000000000";
                when x"1B10" => data <= "0000000000";
                when x"1B11" => data <= "0000000000";
                when x"1B12" => data <= "0000000000";
                when x"1B13" => data <= "0000000000";
                when x"1B14" => data <= "0000000000";
                when x"1B15" => data <= "0000000000";
                when x"1B16" => data <= "0000000000";
                when x"1B17" => data <= "0000000000";
                when x"1B18" => data <= "0000000000";
                when x"1B19" => data <= "0000000000";
                when x"1B1A" => data <= "0000000000";
                when x"1B1B" => data <= "0000000000";
                when x"1B1C" => data <= "0000000000";
                when x"1B1D" => data <= "0000000000";
                when x"1B1E" => data <= "0000000000";
                when x"1B1F" => data <= "0000000000";
                when x"1B20" => data <= "0000000000";
                when x"1B21" => data <= "0000000000";
                when x"1B22" => data <= "0000000000";
                when x"1B23" => data <= "0000000000";
                when x"1B24" => data <= "0000000000";
                when x"1B25" => data <= "0000000000";
                when x"1B26" => data <= "0000000000";
                when x"1B27" => data <= "0000000000";
                when x"1B28" => data <= "0000000000";
                when x"1B29" => data <= "0000000000";
                when x"1B2A" => data <= "0000000000";
                when x"1B2B" => data <= "0000000000";
                when x"1B2C" => data <= "0000000000";
                when x"1B2D" => data <= "0000000000";
                when x"1B2E" => data <= "0000000000";
                when x"1B2F" => data <= "0000000000";
                when x"1B30" => data <= "0000000000";
                when x"1B31" => data <= "0000000000";
                when x"1B32" => data <= "0000000000";
                when x"1B33" => data <= "0000000000";
                when x"1B34" => data <= "0000000000";
                when x"1B35" => data <= "0000000000";
                when x"1B36" => data <= "0000000000";
                when x"1B37" => data <= "0000000000";
                when x"1B38" => data <= "0000000000";
                when x"1B39" => data <= "0000000000";
                when x"1B3A" => data <= "0000000000";
                when x"1B3B" => data <= "0000000000";
                when x"1B3C" => data <= "0000000000";
                when x"1B3D" => data <= "0000000000";
                when x"1B3E" => data <= "0000000000";
                when x"1B3F" => data <= "0000000000";
                when x"1B40" => data <= "0000000000";
                when x"1B41" => data <= "0000000000";
                when x"1B42" => data <= "0000000000";
                when x"1B43" => data <= "0000000000";
                when x"1B44" => data <= "0000000000";
                when x"1B45" => data <= "0000000000";
                when x"1B46" => data <= "0000000000";
                when x"1B47" => data <= "0000000000";
                when x"1B48" => data <= "0000000000";
                when x"1B49" => data <= "0000000000";
                when x"1B4A" => data <= "0000000000";
                when x"1B4B" => data <= "0000000000";
                when x"1B4C" => data <= "0000000000";
                when x"1B4D" => data <= "0000000000";
                when x"1B4E" => data <= "0000000000";
                when x"1B4F" => data <= "0000000000";
                when x"1B50" => data <= "0000000000";
                when x"1B51" => data <= "0000000000";
                when x"1B52" => data <= "0000000000";
                when x"1B53" => data <= "0000000000";
                when x"1B54" => data <= "0000000000";
                when x"1B55" => data <= "0000000000";
                when x"1B56" => data <= "0000000000";
                when x"1B57" => data <= "0000000000";
                when x"1B58" => data <= "0000000000";
                when x"1B59" => data <= "0000000000";
                when x"1B5A" => data <= "0000000000";
                when x"1B5B" => data <= "0000000000";
                when x"1B5C" => data <= "0000000000";
                when x"1B5D" => data <= "0000000000";
                when x"1B5E" => data <= "0000000000";
                when x"1B5F" => data <= "0000000000";
                when x"1B60" => data <= "0000000000";
                when x"1B61" => data <= "0000000000";
                when x"1B62" => data <= "0000000000";
                when x"1B63" => data <= "0000000000";
                when x"1B64" => data <= "0000000000";
                when x"1B65" => data <= "0000000000";
                when x"1B66" => data <= "0000000000";
                when x"1B67" => data <= "0000000000";
                when x"1B68" => data <= "0000000000";
                when x"1B69" => data <= "0000000000";
                when x"1B6A" => data <= "0000000000";
                when x"1B6B" => data <= "0000000000";
                when x"1B6C" => data <= "0000000000";
                when x"1B6D" => data <= "0000000000";
                when x"1B6E" => data <= "0000000000";
                when x"1B6F" => data <= "0000000000";
                when x"1B70" => data <= "0000000000";
                when x"1B71" => data <= "0000000000";
                when x"1B72" => data <= "0000000000";
                when x"1B73" => data <= "0000000000";
                when x"1B74" => data <= "0000000000";
                when x"1B75" => data <= "0000000000";
                when x"1B76" => data <= "0000000000";
                when x"1B77" => data <= "0000000000";
                when x"1B78" => data <= "0000000000";
                when x"1B79" => data <= "0000000000";
                when x"1B7A" => data <= "0000000000";
                when x"1B7B" => data <= "0000000000";
                when x"1B7C" => data <= "0000000000";
                when x"1B7D" => data <= "0000000000";
                when x"1B7E" => data <= "0000000000";
                when x"1B7F" => data <= "0000000000";
                when x"1B80" => data <= "0000000000";
                when x"1B81" => data <= "1010100111";
                when x"1B82" => data <= "0000000000";
                when x"1B83" => data <= "0000000000";
                when x"1B84" => data <= "0000000000";
                when x"1B85" => data <= "0000000000";
                when x"1B86" => data <= "0000000000";
                when x"1B87" => data <= "0000000000";
                when x"1B88" => data <= "0000000000";
                when x"1B89" => data <= "0000000000";
                when x"1B8A" => data <= "0000000000";
                when x"1B8B" => data <= "0000000000";
                when x"1B8C" => data <= "0000000000";
                when x"1B8D" => data <= "0000000000";
                when x"1B8E" => data <= "0000000000";
                when x"1B8F" => data <= "0000000000";
                when x"1B90" => data <= "0000000000";
                when x"1B91" => data <= "0000000000";
                when x"1B92" => data <= "0000000000";
                when x"1B93" => data <= "0000000000";
                when x"1B94" => data <= "0000000000";
                when x"1B95" => data <= "0000000000";
                when x"1B96" => data <= "0000000000";
                when x"1B97" => data <= "0000000000";
                when x"1B98" => data <= "0000000000";
                when x"1B99" => data <= "0000000000";
                when x"1B9A" => data <= "0000000000";
                when x"1B9B" => data <= "0000000000";
                when x"1B9C" => data <= "0000000000";
                when x"1B9D" => data <= "0000000000";
                when x"1B9E" => data <= "0000000000";
                when x"1B9F" => data <= "0000000000";
                when x"1BA0" => data <= "0000000000";
                when x"1BA1" => data <= "0000000000";
                when x"1BA2" => data <= "0000000000";
                when x"1BA3" => data <= "0000000000";
                when x"1BA4" => data <= "0000000000";
                when x"1BA5" => data <= "0000000000";
                when x"1BA6" => data <= "0000000000";
                when x"1BA7" => data <= "0000000000";
                when x"1BA8" => data <= "0000000000";
                when x"1BA9" => data <= "0000000000";
                when x"1BAA" => data <= "0000000000";
                when x"1BAB" => data <= "0000000000";
                when x"1BAC" => data <= "0000000000";
                when x"1BAD" => data <= "0000000000";
                when x"1BAE" => data <= "0000000000";
                when x"1BAF" => data <= "0000000000";
                when x"1BB0" => data <= "0000000000";
                when x"1BB1" => data <= "0000000000";
                when x"1BB2" => data <= "0000000000";
                when x"1BB3" => data <= "0000000000";
                when x"1BB4" => data <= "0000000000";
                when x"1BB5" => data <= "0000000000";
                when x"1BB6" => data <= "0000000000";
                when x"1BB7" => data <= "0000000000";
                when x"1BB8" => data <= "0000000000";
                when x"1BB9" => data <= "0000000000";
                when x"1BBA" => data <= "0000000000";
                when x"1BBB" => data <= "0000000000";
                when x"1BBC" => data <= "0000000000";
                when x"1BBD" => data <= "0000000000";
                when x"1BBE" => data <= "0000000000";
                when x"1BBF" => data <= "0000000000";
                when x"1BC0" => data <= "0000000000";
                when x"1BC1" => data <= "0000000000";
                when x"1BC2" => data <= "0000000000";
                when x"1BC3" => data <= "0000000000";
                when x"1BC4" => data <= "0000000000";
                when x"1BC5" => data <= "0000000000";
                when x"1BC6" => data <= "0000000000";
                when x"1BC7" => data <= "0000000000";
                when x"1BC8" => data <= "0000000000";
                when x"1BC9" => data <= "0000000000";
                when x"1BCA" => data <= "0000000000";
                when x"1BCB" => data <= "0000000000";
                when x"1BCC" => data <= "0000000000";
                when x"1BCD" => data <= "0000000000";
                when x"1BCE" => data <= "0000000000";
                when x"1BCF" => data <= "0000000000";
                when x"1BD0" => data <= "0000000000";
                when x"1BD1" => data <= "0000000000";
                when x"1BD2" => data <= "0000000000";
                when x"1BD3" => data <= "0000000000";
                when x"1BD4" => data <= "0000000000";
                when x"1BD5" => data <= "0000000000";
                when x"1BD6" => data <= "0000000000";
                when x"1BD7" => data <= "0000000000";
                when x"1BD8" => data <= "0000000000";
                when x"1BD9" => data <= "0000000000";
                when x"1BDA" => data <= "0000000000";
                when x"1BDB" => data <= "1011001101";
                when x"1BDC" => data <= "0000000000";
                when x"1BDD" => data <= "0000000000";
                when x"1BDE" => data <= "0000000000";
                when x"1BDF" => data <= "0000000000";
                when x"1BE0" => data <= "0000000000";
                when x"1BE1" => data <= "0000000000";
                when x"1BE2" => data <= "0000000000";
                when x"1BE3" => data <= "0000000000";
                when x"1BE4" => data <= "0000000000";
                when x"1BE5" => data <= "0000000000";
                when x"1BE6" => data <= "0000000000";
                when x"1BE7" => data <= "0000000000";
                when x"1BE8" => data <= "0000000000";
                when x"1BE9" => data <= "0000000000";
                when x"1BEA" => data <= "0000000000";
                when x"1BEB" => data <= "0000000000";
                when x"1BEC" => data <= "0000000000";
                when x"1BED" => data <= "0000000000";
                when x"1BEE" => data <= "0000000000";
                when x"1BEF" => data <= "0000000000";
                when x"1BF0" => data <= "0000000000";
                when x"1BF1" => data <= "0000000000";
                when x"1BF2" => data <= "0000000000";
                when x"1BF3" => data <= "0000000000";
                when x"1BF4" => data <= "0000000000";
                when x"1BF5" => data <= "0000000000";
                when x"1BF6" => data <= "0000000000";
                when x"1BF7" => data <= "0000000000";
                when x"1BF8" => data <= "0000000000";
                when x"1BF9" => data <= "0000000000";
                when x"1BFA" => data <= "0000000000";
                when x"1BFB" => data <= "0000000000";
                when x"1BFC" => data <= "0000000000";
                when x"1BFD" => data <= "0000000000";
                when x"1BFE" => data <= "0000000000";
                when x"1BFF" => data <= "0000000000";
                when x"1C00" => data <= "0000000000";
                when x"1C01" => data <= "0000000000";
                when x"1C02" => data <= "0000000000";
                when x"1C03" => data <= "0000000000";
                when x"1C04" => data <= "0000000000";
                when x"1C05" => data <= "0000000000";
                when x"1C06" => data <= "0000000000";
                when x"1C07" => data <= "0000000000";
                when x"1C08" => data <= "0000000000";
                when x"1C09" => data <= "0000000000";
                when x"1C0A" => data <= "0000000000";
                when x"1C0B" => data <= "0000000000";
                when x"1C0C" => data <= "0000000000";
                when x"1C0D" => data <= "0000000000";
                when x"1C0E" => data <= "0000000000";
                when x"1C0F" => data <= "0000000000";
                when x"1C10" => data <= "0000000000";
                when x"1C11" => data <= "0111110111";
                when x"1C12" => data <= "0000000000";
                when x"1C13" => data <= "0000000000";
                when x"1C14" => data <= "0000000000";
                when x"1C15" => data <= "0111110111";
                when x"1C16" => data <= "0000000000";
                when x"1C17" => data <= "0000000000";
                when x"1C18" => data <= "0000000000";
                when x"1C19" => data <= "0000000000";
                when x"1C1A" => data <= "0000000000";
                when x"1C1B" => data <= "0000000000";
                when x"1C1C" => data <= "0000000000";
                when x"1C1D" => data <= "0000000000";
                when x"1C1E" => data <= "0000000000";
                when x"1C1F" => data <= "0000000000";
                when x"1C20" => data <= "0000000000";
                when x"1C21" => data <= "0000000000";
                when x"1C22" => data <= "0000000000";
                when x"1C23" => data <= "0000000000";
                when x"1C24" => data <= "0000000000";
                when x"1C25" => data <= "0000000000";
                when x"1C26" => data <= "0000000000";
                when x"1C27" => data <= "0000000000";
                when x"1C28" => data <= "0000000000";
                when x"1C29" => data <= "0000000000";
                when x"1C2A" => data <= "0000000000";
                when x"1C2B" => data <= "0000000000";
                when x"1C2C" => data <= "0000000000";
                when x"1C2D" => data <= "0000000000";
                when x"1C2E" => data <= "0000000000";
                when x"1C2F" => data <= "0000000000";
                when x"1C30" => data <= "0000000000";
                when x"1C31" => data <= "0000000000";
                when x"1C32" => data <= "0000000000";
                when x"1C33" => data <= "0000000000";
                when x"1C34" => data <= "0000000000";
                when x"1C35" => data <= "0000000000";
                when x"1C36" => data <= "0000000000";
                when x"1C37" => data <= "0000000000";
                when x"1C38" => data <= "0000000000";
                when x"1C39" => data <= "0000000000";
                when x"1C3A" => data <= "0000000000";
                when x"1C3B" => data <= "0000000000";
                when x"1C3C" => data <= "0000000000";
                when x"1C3D" => data <= "0000000000";
                when x"1C3E" => data <= "0000000000";
                when x"1C3F" => data <= "0000000000";
                when x"1C40" => data <= "0000000000";
                when x"1C41" => data <= "0000000000";
                when x"1C42" => data <= "0000000000";
                when x"1C43" => data <= "0000000000";
                when x"1C44" => data <= "0000000000";
                when x"1C45" => data <= "0000000000";
                when x"1C46" => data <= "0000000000";
                when x"1C47" => data <= "0000000000";
                when x"1C48" => data <= "0000000000";
                when x"1C49" => data <= "0000000000";
                when x"1C4A" => data <= "0000000000";
                when x"1C4B" => data <= "0000000000";
                when x"1C4C" => data <= "0000000000";
                when x"1C4D" => data <= "0000000000";
                when x"1C4E" => data <= "0000000000";
                when x"1C4F" => data <= "0000000000";
                when x"1C50" => data <= "0000000000";
                when x"1C51" => data <= "0000000000";
                when x"1C52" => data <= "0000000000";
                when x"1C53" => data <= "0000000000";
                when x"1C54" => data <= "0000000000";
                when x"1C55" => data <= "0000000000";
                when x"1C56" => data <= "0000000000";
                when x"1C57" => data <= "0000000000";
                when x"1C58" => data <= "0000000000";
                when x"1C59" => data <= "0000000000";
                when x"1C5A" => data <= "0000000000";
                when x"1C5B" => data <= "0000000000";
                when x"1C5C" => data <= "0000000000";
                when x"1C5D" => data <= "0000000000";
                when x"1C5E" => data <= "0000000000";
                when x"1C5F" => data <= "0000000000";
                when x"1C60" => data <= "0000000000";
                when x"1C61" => data <= "0000000000";
                when x"1C62" => data <= "0000000000";
                when x"1C63" => data <= "0000000000";
                when x"1C64" => data <= "0000000000";
                when x"1C65" => data <= "0000000000";
                when x"1C66" => data <= "0000000000";
                when x"1C67" => data <= "0000000000";
                when x"1C68" => data <= "0000000000";
                when x"1C69" => data <= "0000000000";
                when x"1C6A" => data <= "0000000000";
                when x"1C6B" => data <= "0000000000";
                when x"1C6C" => data <= "0000000000";
                when x"1C6D" => data <= "0000000000";
                when x"1C6E" => data <= "0000000000";
                when x"1C6F" => data <= "0000000000";
                when x"1C70" => data <= "0000000000";
                when x"1C71" => data <= "0000000000";
                when x"1C72" => data <= "0000000000";
                when x"1C73" => data <= "0000000000";
                when x"1C74" => data <= "0000000000";
                when x"1C75" => data <= "0000000000";
                when x"1C76" => data <= "0000000000";
                when x"1C77" => data <= "0011100001";
                when x"1C78" => data <= "0000000000";
                when x"1C79" => data <= "0000000000";
                when x"1C7A" => data <= "0000000000";
                when x"1C7B" => data <= "0000000000";
                when x"1C7C" => data <= "0000000000";
                when x"1C7D" => data <= "0000000000";
                when x"1C7E" => data <= "0000000000";
                when x"1C7F" => data <= "0000000000";
                when x"1C80" => data <= "0000000000";
                when x"1C81" => data <= "0000000000";
                when x"1C82" => data <= "0000000000";
                when x"1C83" => data <= "0000000000";
                when x"1C84" => data <= "0000000000";
                when x"1C85" => data <= "0000000000";
                when x"1C86" => data <= "0000000000";
                when x"1C87" => data <= "0000000000";
                when x"1C88" => data <= "0000000000";
                when x"1C89" => data <= "0000000000";
                when x"1C8A" => data <= "0000000000";
                when x"1C8B" => data <= "0000000000";
                when x"1C8C" => data <= "0000000000";
                when x"1C8D" => data <= "0000000000";
                when x"1C8E" => data <= "0000000000";
                when x"1C8F" => data <= "0000000000";
                when x"1C90" => data <= "0000000000";
                when x"1C91" => data <= "0000000000";
                when x"1C92" => data <= "0000000000";
                when x"1C93" => data <= "0000000000";
                when x"1C94" => data <= "0000000000";
                when x"1C95" => data <= "0000000000";
                when x"1C96" => data <= "0000000000";
                when x"1C97" => data <= "0000000000";
                when x"1C98" => data <= "0000000000";
                when x"1C99" => data <= "0000000000";
                when x"1C9A" => data <= "0000000000";
                when x"1C9B" => data <= "0000000000";
                when x"1C9C" => data <= "0000000000";
                when x"1C9D" => data <= "0000000000";
                when x"1C9E" => data <= "0000000000";
                when x"1C9F" => data <= "0000000000";
                when x"1CA0" => data <= "0000000000";
                when x"1CA1" => data <= "0000000000";
                when x"1CA2" => data <= "0000000000";
                when x"1CA3" => data <= "0000000000";
                when x"1CA4" => data <= "0000000000";
                when x"1CA5" => data <= "0000000000";
                when x"1CA6" => data <= "0000000000";
                when x"1CA7" => data <= "0000000000";
                when x"1CA8" => data <= "0000000000";
                when x"1CA9" => data <= "0000000000";
                when x"1CAA" => data <= "0000000000";
                when x"1CAB" => data <= "0000000000";
                when x"1CAC" => data <= "0000000000";
                when x"1CAD" => data <= "0000000000";
                when x"1CAE" => data <= "0000000000";
                when x"1CAF" => data <= "0000000000";
                when x"1CB0" => data <= "0000000000";
                when x"1CB1" => data <= "0000000000";
                when x"1CB2" => data <= "0000000000";
                when x"1CB3" => data <= "0000000000";
                when x"1CB4" => data <= "0000000000";
                when x"1CB5" => data <= "0000000000";
                when x"1CB6" => data <= "0000000000";
                when x"1CB7" => data <= "0000000000";
                when x"1CB8" => data <= "0000000000";
                when x"1CB9" => data <= "0000000000";
                when x"1CBA" => data <= "0000000000";
                when x"1CBB" => data <= "0000000000";
                when x"1CBC" => data <= "0000000000";
                when x"1CBD" => data <= "0000000000";
                when x"1CBE" => data <= "0000000000";
                when x"1CBF" => data <= "0000000000";
                when x"1CC0" => data <= "0000000000";
                when x"1CC1" => data <= "0000000000";
                when x"1CC2" => data <= "0000000000";
                when x"1CC3" => data <= "0000000000";
                when x"1CC4" => data <= "0000000000";
                when x"1CC5" => data <= "0000000000";
                when x"1CC6" => data <= "0000000000";
                when x"1CC7" => data <= "0000000000";
                when x"1CC8" => data <= "0000000000";
                when x"1CC9" => data <= "0000000000";
                when x"1CCA" => data <= "0000000000";
                when x"1CCB" => data <= "0000000000";
                when x"1CCC" => data <= "0000000000";
                when x"1CCD" => data <= "0000000000";
                when x"1CCE" => data <= "0000000000";
                when x"1CCF" => data <= "0000000000";
                when x"1CD0" => data <= "0000000000";
                when x"1CD1" => data <= "0000000000";
                when x"1CD2" => data <= "0000000000";
                when x"1CD3" => data <= "0000000000";
                when x"1CD4" => data <= "0000000000";
                when x"1CD5" => data <= "0000000000";
                when x"1CD6" => data <= "0000000000";
                when x"1CD7" => data <= "0000000000";
                when x"1CD8" => data <= "0000000000";
                when x"1CD9" => data <= "0000000000";
                when x"1CDA" => data <= "0000000000";
                when x"1CDB" => data <= "0000000000";
                when x"1CDC" => data <= "0000000000";
                when x"1CDD" => data <= "0000000000";
                when x"1CDE" => data <= "0000000000";
                when x"1CDF" => data <= "0000000000";
                when x"1CE0" => data <= "0000000000";
                when x"1CE1" => data <= "0000000000";
                when x"1CE2" => data <= "0000000000";
                when x"1CE3" => data <= "0000000000";
                when x"1CE4" => data <= "0000000000";
                when x"1CE5" => data <= "0000000000";
                when x"1CE6" => data <= "0000000000";
                when x"1CE7" => data <= "0000000000";
                when x"1CE8" => data <= "0000000000";
                when x"1CE9" => data <= "0000000000";
                when x"1CEA" => data <= "0000000000";
                when x"1CEB" => data <= "0000000000";
                when x"1CEC" => data <= "0000000000";
                when x"1CED" => data <= "0000000000";
                when x"1CEE" => data <= "0000000000";
                when x"1CEF" => data <= "0000000000";
                when x"1CF0" => data <= "0000000000";
                when x"1CF1" => data <= "0000000000";
                when x"1CF2" => data <= "0000000000";
                when x"1CF3" => data <= "0000000000";
                when x"1CF4" => data <= "0000000000";
                when x"1CF5" => data <= "0000000000";
                when x"1CF6" => data <= "0000000000";
                when x"1CF7" => data <= "0000000000";
                when x"1CF8" => data <= "0000000000";
                when x"1CF9" => data <= "0000000000";
                when x"1CFA" => data <= "0000000000";
                when x"1CFB" => data <= "0000000000";
                when x"1CFC" => data <= "0000000000";
                when x"1CFD" => data <= "0000000000";
                when x"1CFE" => data <= "0000000000";
                when x"1CFF" => data <= "0000000000";
                when x"1D00" => data <= "0000000000";
                when x"1D01" => data <= "0000000000";
                when x"1D02" => data <= "0000000000";
                when x"1D03" => data <= "0000000000";
                when x"1D04" => data <= "0000000000";
                when x"1D05" => data <= "0000000000";
                when x"1D06" => data <= "0000000000";
                when x"1D07" => data <= "0000000000";
                when x"1D08" => data <= "0000000000";
                when x"1D09" => data <= "0000000000";
                when x"1D0A" => data <= "0000000000";
                when x"1D0B" => data <= "0000000000";
                when x"1D0C" => data <= "0000000000";
                when x"1D0D" => data <= "0000000000";
                when x"1D0E" => data <= "0000000000";
                when x"1D0F" => data <= "0000000000";
                when x"1D10" => data <= "1000101100";
                when x"1D11" => data <= "0000000000";
                when x"1D12" => data <= "0000000000";
                when x"1D13" => data <= "0000000000";
                when x"1D14" => data <= "0000000000";
                when x"1D15" => data <= "0000000000";
                when x"1D16" => data <= "0000000000";
                when x"1D17" => data <= "0000000000";
                when x"1D18" => data <= "0000000000";
                when x"1D19" => data <= "0000000000";
                when x"1D1A" => data <= "0000000000";
                when x"1D1B" => data <= "0000000000";
                when x"1D1C" => data <= "0000000000";
                when x"1D1D" => data <= "0000000000";
                when x"1D1E" => data <= "0000000000";
                when x"1D1F" => data <= "0000000000";
                when x"1D20" => data <= "0000000000";
                when x"1D21" => data <= "0000000000";
                when x"1D22" => data <= "0000000000";
                when x"1D23" => data <= "0000000000";
                when x"1D24" => data <= "0000000000";
                when x"1D25" => data <= "0000000000";
                when x"1D26" => data <= "0000000000";
                when x"1D27" => data <= "0000000000";
                when x"1D28" => data <= "0000000000";
                when x"1D29" => data <= "0000000000";
                when x"1D2A" => data <= "0000000000";
                when x"1D2B" => data <= "0000000000";
                when x"1D2C" => data <= "0000000000";
                when x"1D2D" => data <= "0000000000";
                when x"1D2E" => data <= "0000000000";
                when x"1D2F" => data <= "0000000000";
                when x"1D30" => data <= "0000000000";
                when x"1D31" => data <= "0000000000";
                when x"1D32" => data <= "0000000000";
                when x"1D33" => data <= "0000000000";
                when x"1D34" => data <= "0000000000";
                when x"1D35" => data <= "0000000000";
                when x"1D36" => data <= "1111011011";
                when x"1D37" => data <= "0000000000";
                when x"1D38" => data <= "0000000000";
                when x"1D39" => data <= "0000000000";
                when x"1D3A" => data <= "0000000000";
                when x"1D3B" => data <= "0000000000";
                when x"1D3C" => data <= "0000000000";
                when x"1D3D" => data <= "0000000000";
                when x"1D3E" => data <= "0000000000";
                when x"1D3F" => data <= "0000000000";
                when x"1D40" => data <= "0000000000";
                when x"1D41" => data <= "0000000000";
                when x"1D42" => data <= "0000000000";
                when x"1D43" => data <= "0000000000";
                when x"1D44" => data <= "0000000000";
                when x"1D45" => data <= "0000000000";
                when x"1D46" => data <= "0000000000";
                when x"1D47" => data <= "0000000000";
                when x"1D48" => data <= "0000000000";
                when x"1D49" => data <= "0000000000";
                when x"1D4A" => data <= "0000000000";
                when x"1D4B" => data <= "0000000000";
                when x"1D4C" => data <= "0000000000";
                when x"1D4D" => data <= "0000000000";
                when x"1D4E" => data <= "0000000000";
                when x"1D4F" => data <= "0000000000";
                when x"1D50" => data <= "0000000000";
                when x"1D51" => data <= "0000000000";
                when x"1D52" => data <= "0000000000";
                when x"1D53" => data <= "0000000000";
                when x"1D54" => data <= "0000000000";
                when x"1D55" => data <= "0000000000";
                when x"1D56" => data <= "1111011011";
                when x"1D57" => data <= "0000000000";
                when x"1D58" => data <= "0000000000";
                when x"1D59" => data <= "0000000000";
                when x"1D5A" => data <= "0000000000";
                when x"1D5B" => data <= "0000000000";
                when x"1D5C" => data <= "0000000000";
                when x"1D5D" => data <= "0000000000";
                when x"1D5E" => data <= "0000000000";
                when x"1D5F" => data <= "0000000000";
                when x"1D60" => data <= "0000000000";
                when x"1D61" => data <= "0000000000";
                when x"1D62" => data <= "0000000000";
                when x"1D63" => data <= "0000000000";
                when x"1D64" => data <= "0000000000";
                when x"1D65" => data <= "0000000000";
                when x"1D66" => data <= "0000000000";
                when x"1D67" => data <= "0000000000";
                when x"1D68" => data <= "0000000000";
                when x"1D69" => data <= "1111011011";
                when x"1D6A" => data <= "0000000000";
                when x"1D6B" => data <= "0000000000";
                when x"1D6C" => data <= "0000000000";
                when x"1D6D" => data <= "0000000000";
                when x"1D6E" => data <= "0000000000";
                when x"1D6F" => data <= "0000000000";
                when x"1D70" => data <= "0000000000";
                when x"1D71" => data <= "0000000000";
                when x"1D72" => data <= "0000000000";
                when x"1D73" => data <= "0000000000";
                when x"1D74" => data <= "0000000000";
                when x"1D75" => data <= "0000000000";
                when x"1D76" => data <= "0000000000";
                when x"1D77" => data <= "0000000000";
                when x"1D78" => data <= "0000000000";
                when x"1D79" => data <= "0000000000";
                when x"1D7A" => data <= "0000000000";
                when x"1D7B" => data <= "0000000000";
                when x"1D7C" => data <= "0000000000";
                when x"1D7D" => data <= "0100100011";
                when x"1D7E" => data <= "0000000000";
                when x"1D7F" => data <= "0000000000";
                when x"1D80" => data <= "0000000000";
                when x"1D81" => data <= "0000000000";
                when x"1D82" => data <= "0000000000";
                when x"1D83" => data <= "0000000000";
                when x"1D84" => data <= "0000000000";
                when x"1D85" => data <= "0000000000";
                when x"1D86" => data <= "0000000000";
                when x"1D87" => data <= "0000000000";
                when x"1D88" => data <= "0000000000";
                when x"1D89" => data <= "0000000000";
                when x"1D8A" => data <= "0000000000";
                when x"1D8B" => data <= "0000000000";
                when x"1D8C" => data <= "0000000000";
                when x"1D8D" => data <= "0000000000";
                when x"1D8E" => data <= "0000000000";
                when x"1D8F" => data <= "0000000000";
                when x"1D90" => data <= "0000000000";
                when x"1D91" => data <= "0000000000";
                when x"1D92" => data <= "0000000000";
                when x"1D93" => data <= "0000000000";
                when x"1D94" => data <= "0000000000";
                when x"1D95" => data <= "0000000000";
                when x"1D96" => data <= "0000000000";
                when x"1D97" => data <= "0000000000";
                when x"1D98" => data <= "0000000000";
                when x"1D99" => data <= "0000000000";
                when x"1D9A" => data <= "0000000000";
                when x"1D9B" => data <= "0000000000";
                when x"1D9C" => data <= "0000000000";
                when x"1D9D" => data <= "0000000000";
                when x"1D9E" => data <= "0000000000";
                when x"1D9F" => data <= "0000000000";
                when x"1DA0" => data <= "0000000000";
                when x"1DA1" => data <= "0000000000";
                when x"1DA2" => data <= "0000000000";
                when x"1DA3" => data <= "0000000000";
                when x"1DA4" => data <= "0000000000";
                when x"1DA5" => data <= "0000000000";
                when x"1DA6" => data <= "0000000000";
                when x"1DA7" => data <= "0000000000";
                when x"1DA8" => data <= "0000000000";
                when x"1DA9" => data <= "0000000000";
                when x"1DAA" => data <= "0000000000";
                when x"1DAB" => data <= "0000000000";
                when x"1DAC" => data <= "0000000000";
                when x"1DAD" => data <= "0000000000";
                when x"1DAE" => data <= "0000000000";
                when x"1DAF" => data <= "0000000000";
                when x"1DB0" => data <= "0000000000";
                when x"1DB1" => data <= "0000000000";
                when x"1DB2" => data <= "0000000000";
                when x"1DB3" => data <= "0000000000";
                when x"1DB4" => data <= "0000000000";
                when x"1DB5" => data <= "0000000000";
                when x"1DB6" => data <= "0000000000";
                when x"1DB7" => data <= "0000000000";
                when x"1DB8" => data <= "0000000000";
                when x"1DB9" => data <= "0000000000";
                when x"1DBA" => data <= "0000000000";
                when x"1DBB" => data <= "0000000000";
                when x"1DBC" => data <= "0000000000";
                when x"1DBD" => data <= "0000000000";
                when x"1DBE" => data <= "0000000000";
                when x"1DBF" => data <= "0000000000";
                when x"1DC0" => data <= "0000000000";
                when x"1DC1" => data <= "0000000000";
                when x"1DC2" => data <= "0000000000";
                when x"1DC3" => data <= "0000000000";
                when x"1DC4" => data <= "0000000000";
                when x"1DC5" => data <= "0000000000";
                when x"1DC6" => data <= "0000000000";
                when x"1DC7" => data <= "0000000000";
                when x"1DC8" => data <= "0000000000";
                when x"1DC9" => data <= "0000000000";
                when x"1DCA" => data <= "0000000000";
                when x"1DCB" => data <= "0000000000";
                when x"1DCC" => data <= "0000000000";
                when x"1DCD" => data <= "0000000000";
                when x"1DCE" => data <= "1011001101";
                when x"1DCF" => data <= "0000000000";
                when x"1DD0" => data <= "0000000000";
                when x"1DD1" => data <= "0000000000";
                when x"1DD2" => data <= "0000000000";
                when x"1DD3" => data <= "0000000000";
                when x"1DD4" => data <= "0000000000";
                when x"1DD5" => data <= "0000000000";
                when x"1DD6" => data <= "0000000000";
                when x"1DD7" => data <= "0000000000";
                when x"1DD8" => data <= "0000000000";
                when x"1DD9" => data <= "0000000000";
                when x"1DDA" => data <= "0000000000";
                when x"1DDB" => data <= "0000000000";
                when x"1DDC" => data <= "0000000000";
                when x"1DDD" => data <= "0000000000";
                when x"1DDE" => data <= "0000000000";
                when x"1DDF" => data <= "0000000000";
                when x"1DE0" => data <= "0000000000";
                when x"1DE1" => data <= "0000000000";
                when x"1DE2" => data <= "0000000000";
                when x"1DE3" => data <= "0000000000";
                when x"1DE4" => data <= "0000000000";
                when x"1DE5" => data <= "0000000000";
                when x"1DE6" => data <= "0000000000";
                when x"1DE7" => data <= "0000000000";
                when x"1DE8" => data <= "0000000000";
                when x"1DE9" => data <= "0000000000";
                when x"1DEA" => data <= "0000000000";
                when x"1DEB" => data <= "0000000000";
                when x"1DEC" => data <= "0000000000";
                when x"1DED" => data <= "0000000000";
                when x"1DEE" => data <= "0000000000";
                when x"1DEF" => data <= "0000000000";
                when x"1DF0" => data <= "0000000000";
                when x"1DF1" => data <= "0000000000";
                when x"1DF2" => data <= "0000000000";
                when x"1DF3" => data <= "0000000000";
                when x"1DF4" => data <= "0000000000";
                when x"1DF5" => data <= "0000000000";
                when x"1DF6" => data <= "0000000000";
                when x"1DF7" => data <= "0000000000";
                when x"1DF8" => data <= "0000000000";
                when x"1DF9" => data <= "0000000000";
                when x"1DFA" => data <= "0000000000";
                when x"1DFB" => data <= "0000000000";
                when x"1DFC" => data <= "0000000000";
                when x"1DFD" => data <= "0000000000";
                when x"1DFE" => data <= "0000000000";
                when x"1DFF" => data <= "0000000000";
                when x"1E00" => data <= "0000000000";
                when x"1E01" => data <= "0000000000";
                when x"1E02" => data <= "0000000000";
                when x"1E03" => data <= "0000000000";
                when x"1E04" => data <= "0000000000";
                when x"1E05" => data <= "0000000000";
                when x"1E06" => data <= "0000000000";
                when x"1E07" => data <= "0000000000";
                when x"1E08" => data <= "0000000000";
                when x"1E09" => data <= "0000000000";
                when x"1E0A" => data <= "0000000000";
                when x"1E0B" => data <= "0000000000";
                when x"1E0C" => data <= "0000000000";
                when x"1E0D" => data <= "0000000000";
                when x"1E0E" => data <= "0000000000";
                when x"1E0F" => data <= "0000000000";
                when x"1E10" => data <= "0000000000";
                when x"1E11" => data <= "0000000000";
                when x"1E12" => data <= "0111110111";
                when x"1E13" => data <= "0000000000";
                when x"1E14" => data <= "0000000000";
                when x"1E15" => data <= "0000000000";
                when x"1E16" => data <= "0000000000";
                when x"1E17" => data <= "0000000000";
                when x"1E18" => data <= "0000000000";
                when x"1E19" => data <= "0000000000";
                when x"1E1A" => data <= "0000000000";
                when x"1E1B" => data <= "0000000000";
                when x"1E1C" => data <= "0000000000";
                when x"1E1D" => data <= "0000000000";
                when x"1E1E" => data <= "0000000000";
                when x"1E1F" => data <= "0000000000";
                when x"1E20" => data <= "0000000000";
                when x"1E21" => data <= "0000000000";
                when x"1E22" => data <= "0000000000";
                when x"1E23" => data <= "0000000000";
                when x"1E24" => data <= "0000000000";
                when x"1E25" => data <= "0000000000";
                when x"1E26" => data <= "0000000000";
                when x"1E27" => data <= "0000000000";
                when x"1E28" => data <= "0000000000";
                when x"1E29" => data <= "0000000000";
                when x"1E2A" => data <= "0000000000";
                when x"1E2B" => data <= "0000000000";
                when x"1E2C" => data <= "0000000000";
                when x"1E2D" => data <= "0000000000";
                when x"1E2E" => data <= "0000000000";
                when x"1E2F" => data <= "0000000000";
                when x"1E30" => data <= "0000000000";
                when x"1E31" => data <= "0000000000";
                when x"1E32" => data <= "0000000000";
                when x"1E33" => data <= "0000000000";
                when x"1E34" => data <= "0000000000";
                when x"1E35" => data <= "0000000000";
                when x"1E36" => data <= "0000000000";
                when x"1E37" => data <= "0000000000";
                when x"1E38" => data <= "0000000000";
                when x"1E39" => data <= "0000000000";
                when x"1E3A" => data <= "0000000000";
                when x"1E3B" => data <= "0000000000";
                when x"1E3C" => data <= "0000000000";
                when x"1E3D" => data <= "0000000000";
                when x"1E3E" => data <= "0000000000";
                when x"1E3F" => data <= "0000000000";
                when x"1E40" => data <= "0000000000";
                when x"1E41" => data <= "0000000000";
                when x"1E42" => data <= "0000000000";
                when x"1E43" => data <= "0000000000";
                when x"1E44" => data <= "0000000000";
                when x"1E45" => data <= "0000000000";
                when x"1E46" => data <= "0000000000";
                when x"1E47" => data <= "0000000000";
                when x"1E48" => data <= "0000000000";
                when x"1E49" => data <= "0000000000";
                when x"1E4A" => data <= "1101010000";
                when x"1E4B" => data <= "0000000000";
                when x"1E4C" => data <= "0000000000";
                when x"1E4D" => data <= "0000000000";
                when x"1E4E" => data <= "0000000000";
                when x"1E4F" => data <= "0000000000";
                when x"1E50" => data <= "0000000000";
                when x"1E51" => data <= "0000000000";
                when x"1E52" => data <= "0000000000";
                when x"1E53" => data <= "0000000000";
                when x"1E54" => data <= "0000000000";
                when x"1E55" => data <= "0000000000";
                when x"1E56" => data <= "0000000000";
                when x"1E57" => data <= "0000000000";
                when x"1E58" => data <= "0000000000";
                when x"1E59" => data <= "0000000000";
                when x"1E5A" => data <= "0000000000";
                when x"1E5B" => data <= "0000000000";
                when x"1E5C" => data <= "0000000000";
                when x"1E5D" => data <= "0000000000";
                when x"1E5E" => data <= "0000000000";
                when x"1E5F" => data <= "0000000000";
                when x"1E60" => data <= "0000000000";
                when x"1E61" => data <= "0000000000";
                when x"1E62" => data <= "0000000000";
                when x"1E63" => data <= "0000000000";
                when x"1E64" => data <= "0000000000";
                when x"1E65" => data <= "0000000000";
                when x"1E66" => data <= "0000000000";
                when x"1E67" => data <= "0000000000";
                when x"1E68" => data <= "0000000000";
                when x"1E69" => data <= "0000000000";
                when x"1E6A" => data <= "0000000000";
                when x"1E6B" => data <= "0000000000";
                when x"1E6C" => data <= "0000000000";
                when x"1E6D" => data <= "0000000000";
                when x"1E6E" => data <= "0000000000";
                when x"1E6F" => data <= "0000000000";
                when x"1E70" => data <= "0000000000";
                when x"1E71" => data <= "0000000000";
                when x"1E72" => data <= "0000000000";
                when x"1E73" => data <= "0000000000";
                when x"1E74" => data <= "0000000000";
                when x"1E75" => data <= "0000000000";
                when x"1E76" => data <= "0000000000";
                when x"1E77" => data <= "0000000000";
                when x"1E78" => data <= "0000000000";
                when x"1E79" => data <= "0000000000";
                when x"1E7A" => data <= "0000000000";
                when x"1E7B" => data <= "0000000000";
                when x"1E7C" => data <= "0000000000";
                when x"1E7D" => data <= "0000000000";
                when x"1E7E" => data <= "0000000000";
                when x"1E7F" => data <= "0000000000";
                when x"1E80" => data <= "0000000000";
                when x"1E81" => data <= "0000000000";
                when x"1E82" => data <= "0000000000";
                when x"1E83" => data <= "0000000000";
                when x"1E84" => data <= "0000000000";
                when x"1E85" => data <= "0000000000";
                when x"1E86" => data <= "0000000000";
                when x"1E87" => data <= "0000000000";
                when x"1E88" => data <= "0000000000";
                when x"1E89" => data <= "0000000000";
                when x"1E8A" => data <= "0000000000";
                when x"1E8B" => data <= "0000000000";
                when x"1E8C" => data <= "0000000000";
                when x"1E8D" => data <= "0000000000";
                when x"1E8E" => data <= "0000000000";
                when x"1E8F" => data <= "0000000000";
                when x"1E90" => data <= "0000000000";
                when x"1E91" => data <= "0000000000";
                when x"1E92" => data <= "0000000000";
                when x"1E93" => data <= "0000000000";
                when x"1E94" => data <= "0000000000";
                when x"1E95" => data <= "0000000000";
                when x"1E96" => data <= "0000000000";
                when x"1E97" => data <= "0000000000";
                when x"1E98" => data <= "0000000000";
                when x"1E99" => data <= "0000000000";
                when x"1E9A" => data <= "0000000000";
                when x"1E9B" => data <= "0000000000";
                when x"1E9C" => data <= "0000000000";
                when x"1E9D" => data <= "0000000000";
                when x"1E9E" => data <= "0000000000";
                when x"1E9F" => data <= "0000000000";
                when x"1EA0" => data <= "0000000000";
                when x"1EA1" => data <= "0000000000";
                when x"1EA2" => data <= "0000000000";
                when x"1EA3" => data <= "0000000000";
                when x"1EA4" => data <= "0000000000";
                when x"1EA5" => data <= "0000000000";
                when x"1EA6" => data <= "0000000000";
                when x"1EA7" => data <= "0000000000";
                when x"1EA8" => data <= "0000000000";
                when x"1EA9" => data <= "0000000000";
                when x"1EAA" => data <= "0000000000";
                when x"1EAB" => data <= "0000000000";
                when x"1EAC" => data <= "0000000000";
                when x"1EAD" => data <= "0111110111";
                when x"1EAE" => data <= "0000000000";
                when x"1EAF" => data <= "0000000000";
                when x"1EB0" => data <= "0000000000";
                when x"1EB1" => data <= "0000000000";
                when x"1EB2" => data <= "0000000000";
                when x"1EB3" => data <= "0000000000";
                when x"1EB4" => data <= "0000000000";
                when x"1EB5" => data <= "0000000000";
                when x"1EB6" => data <= "0000000000";
                when x"1EB7" => data <= "0000000000";
                when x"1EB8" => data <= "0000000000";
                when x"1EB9" => data <= "0000000000";
                when x"1EBA" => data <= "0000000000";
                when x"1EBB" => data <= "0000000000";
                when x"1EBC" => data <= "0000000000";
                when x"1EBD" => data <= "0000000000";
                when x"1EBE" => data <= "0000000000";
                when x"1EBF" => data <= "0000000000";
                when x"1EC0" => data <= "0000000000";
                when x"1EC1" => data <= "0000000000";
                when x"1EC2" => data <= "0000000000";
                when x"1EC3" => data <= "0000000000";
                when x"1EC4" => data <= "0000000000";
                when x"1EC5" => data <= "0000000000";
                when x"1EC6" => data <= "0000000000";
                when x"1EC7" => data <= "0000000000";
                when x"1EC8" => data <= "0000000000";
                when x"1EC9" => data <= "0000000000";
                when x"1ECA" => data <= "0000000000";
                when x"1ECB" => data <= "0000000000";
                when x"1ECC" => data <= "0000000000";
                when x"1ECD" => data <= "0000000000";
                when x"1ECE" => data <= "0000000000";
                when x"1ECF" => data <= "0000000000";
                when x"1ED0" => data <= "0000000000";
                when x"1ED1" => data <= "0000000000";
                when x"1ED2" => data <= "0000000000";
                when x"1ED3" => data <= "0000000000";
                when x"1ED4" => data <= "0000000000";
                when x"1ED5" => data <= "0000000000";
                when x"1ED6" => data <= "0000000000";
                when x"1ED7" => data <= "0000000000";
                when x"1ED8" => data <= "0000000000";
                when x"1ED9" => data <= "0000000000";
                when x"1EDA" => data <= "0000000000";
                when x"1EDB" => data <= "0000000000";
                when x"1EDC" => data <= "0000000000";
                when x"1EDD" => data <= "0000000000";
                when x"1EDE" => data <= "0000000000";
                when x"1EDF" => data <= "0000000000";
                when x"1EE0" => data <= "0000000000";
                when x"1EE1" => data <= "0000000000";
                when x"1EE2" => data <= "0000000000";
                when x"1EE3" => data <= "0000000000";
                when x"1EE4" => data <= "0000000000";
                when x"1EE5" => data <= "0000000000";
                when x"1EE6" => data <= "0000000000";
                when x"1EE7" => data <= "0000000000";
                when x"1EE8" => data <= "0000000000";
                when x"1EE9" => data <= "0000000000";
                when x"1EEA" => data <= "0000000000";
                when x"1EEB" => data <= "0000000000";
                when x"1EEC" => data <= "0000000000";
                when x"1EED" => data <= "0000000000";
                when x"1EEE" => data <= "0000000000";
                when x"1EEF" => data <= "0000000000";
                when x"1EF0" => data <= "0000000000";
                when x"1EF1" => data <= "0000000000";
                when x"1EF2" => data <= "0000000000";
                when x"1EF3" => data <= "0000000000";
                when x"1EF4" => data <= "0000000000";
                when x"1EF5" => data <= "0000000000";
                when x"1EF6" => data <= "0000000000";
                when x"1EF7" => data <= "0000000000";
                when x"1EF8" => data <= "0000000000";
                when x"1EF9" => data <= "0000000000";
                when x"1EFA" => data <= "0000000000";
                when x"1EFB" => data <= "0000000000";
                when x"1EFC" => data <= "0000000000";
                when x"1EFD" => data <= "0000000000";
                when x"1EFE" => data <= "0000000000";
                when x"1EFF" => data <= "0000000000";
                when x"1F00" => data <= "0000000000";
                when x"1F01" => data <= "0000000000";
                when x"1F02" => data <= "0000000000";
                when x"1F03" => data <= "0000000000";
                when x"1F04" => data <= "0000000000";
                when x"1F05" => data <= "0000000000";
                when x"1F06" => data <= "0000000000";
                when x"1F07" => data <= "0000000000";
                when x"1F08" => data <= "0000000000";
                when x"1F09" => data <= "0000000000";
                when x"1F0A" => data <= "0000000000";
                when x"1F0B" => data <= "0000000000";
                when x"1F0C" => data <= "0000000000";
                when x"1F0D" => data <= "0000000000";
                when x"1F0E" => data <= "0000000000";
                when x"1F0F" => data <= "0000000000";
                when x"1F10" => data <= "0000000000";
                when x"1F11" => data <= "0000000000";
                when x"1F12" => data <= "0000000000";
                when x"1F13" => data <= "0000000000";
                when x"1F14" => data <= "0000000000";
                when x"1F15" => data <= "0000000000";
                when x"1F16" => data <= "0000000000";
                when x"1F17" => data <= "0000000000";
                when x"1F18" => data <= "0000000000";
                when x"1F19" => data <= "0000000000";
                when x"1F1A" => data <= "0000000000";
                when x"1F1B" => data <= "0000000000";
                when x"1F1C" => data <= "0000000000";
                when x"1F1D" => data <= "0000000000";
                when x"1F1E" => data <= "0000000000";
                when x"1F1F" => data <= "0000000000";
                when x"1F20" => data <= "0000000000";
                when x"1F21" => data <= "0000000000";
                when x"1F22" => data <= "0000000000";
                when x"1F23" => data <= "0000000000";
                when x"1F24" => data <= "0000000000";
                when x"1F25" => data <= "0000000000";
                when x"1F26" => data <= "0000000000";
                when x"1F27" => data <= "0000000000";
                when x"1F28" => data <= "0000000000";
                when x"1F29" => data <= "0000000000";
                when x"1F2A" => data <= "0000000000";
                when x"1F2B" => data <= "0000000000";
                when x"1F2C" => data <= "0000000000";
                when x"1F2D" => data <= "0000000000";
                when x"1F2E" => data <= "0000000000";
                when x"1F2F" => data <= "0000000000";
                when x"1F30" => data <= "0000000000";
                when x"1F31" => data <= "0000000000";
                when x"1F32" => data <= "0000000000";
                when x"1F33" => data <= "0000000000";
                when x"1F34" => data <= "0000000000";
                when x"1F35" => data <= "0000000000";
                when x"1F36" => data <= "0000000000";
                when x"1F37" => data <= "0000000000";
                when x"1F38" => data <= "0000000000";
                when x"1F39" => data <= "0000000000";
                when x"1F3A" => data <= "0000000000";
                when x"1F3B" => data <= "0000000000";
                when x"1F3C" => data <= "0000000000";
                when x"1F3D" => data <= "0000000000";
                when x"1F3E" => data <= "0000000000";
                when x"1F3F" => data <= "0000000000";
                when x"1F40" => data <= "0000000000";
                when x"1F41" => data <= "0000000000";
                when x"1F42" => data <= "0000000000";
                when x"1F43" => data <= "0000000000";
                when x"1F44" => data <= "0000000000";
                when x"1F45" => data <= "0000000000";
                when x"1F46" => data <= "0000000000";
                when x"1F47" => data <= "0000000000";
                when x"1F48" => data <= "0000000000";
                when x"1F49" => data <= "0000000000";
                when x"1F4A" => data <= "0000000000";
                when x"1F4B" => data <= "0000000000";
                when x"1F4C" => data <= "0000000000";
                when x"1F4D" => data <= "0000000000";
                when x"1F4E" => data <= "0000000000";
                when x"1F4F" => data <= "0000000000";
                when x"1F50" => data <= "0000000000";
                when x"1F51" => data <= "0000000000";
                when x"1F52" => data <= "0000000000";
                when x"1F53" => data <= "0000000000";
                when x"1F54" => data <= "0000000000";
                when x"1F55" => data <= "0000000000";
                when x"1F56" => data <= "0000000000";
                when x"1F57" => data <= "0000000000";
                when x"1F58" => data <= "0000000000";
                when x"1F59" => data <= "0000000000";
                when x"1F5A" => data <= "0000000000";
                when x"1F5B" => data <= "0000000000";
                when x"1F5C" => data <= "0000000000";
                when x"1F5D" => data <= "0000000000";
                when x"1F5E" => data <= "0000000000";
                when x"1F5F" => data <= "0000000000";
                when x"1F60" => data <= "0000000000";
                when x"1F61" => data <= "0000000000";
                when x"1F62" => data <= "0000000000";
                when x"1F63" => data <= "0000000000";
                when x"1F64" => data <= "0000000000";
                when x"1F65" => data <= "0000000000";
                when x"1F66" => data <= "0000000000";
                when x"1F67" => data <= "0000000000";
                when x"1F68" => data <= "0111000010";
                when x"1F69" => data <= "0000000000";
                when x"1F6A" => data <= "0000000000";
                when x"1F6B" => data <= "0000000000";
                when x"1F6C" => data <= "0000000000";
                when x"1F6D" => data <= "0000000000";
                when x"1F6E" => data <= "0000000000";
                when x"1F6F" => data <= "0000000000";
                when x"1F70" => data <= "0000000000";
                when x"1F71" => data <= "0000000000";
                when x"1F72" => data <= "0000000000";
                when x"1F73" => data <= "0000000000";
                when x"1F74" => data <= "0000000000";
                when x"1F75" => data <= "0000000000";
                when x"1F76" => data <= "0000000000";
                when x"1F77" => data <= "0000000000";
                when x"1F78" => data <= "0000000000";
                when x"1F79" => data <= "0000000000";
                when x"1F7A" => data <= "0000000000";
                when x"1F7B" => data <= "0000000000";
                when x"1F7C" => data <= "0000000000";
                when x"1F7D" => data <= "0000000000";
                when x"1F7E" => data <= "0000000000";
                when x"1F7F" => data <= "0000000000";
                when x"1F80" => data <= "0000000000";
                when x"1F81" => data <= "0000000000";
                when x"1F82" => data <= "0000000000";
                when x"1F83" => data <= "0000000000";
                when x"1F84" => data <= "0000000000";
                when x"1F85" => data <= "0000000000";
                when x"1F86" => data <= "0000000000";
                when x"1F87" => data <= "0000000000";
                when x"1F88" => data <= "0000000000";
                when x"1F89" => data <= "0000000000";
                when x"1F8A" => data <= "0000000000";
                when x"1F8B" => data <= "0000000000";
                when x"1F8C" => data <= "0000000000";
                when x"1F8D" => data <= "0000000000";
                when x"1F8E" => data <= "0000000000";
                when x"1F8F" => data <= "0000000000";
                when x"1F90" => data <= "0111110111";
                when x"1F91" => data <= "0000000000";
                when x"1F92" => data <= "0000000000";
                when x"1F93" => data <= "0000000000";
                when x"1F94" => data <= "0000000000";
                when x"1F95" => data <= "0000000000";
                when x"1F96" => data <= "0000000000";
                when x"1F97" => data <= "0000000000";
                when x"1F98" => data <= "0000000000";
                when x"1F99" => data <= "0000000000";
                when x"1F9A" => data <= "0000000000";
                when x"1F9B" => data <= "0000000000";
                when x"1F9C" => data <= "0000000000";
                when x"1F9D" => data <= "0000000000";
                when x"1F9E" => data <= "0000000000";
                when x"1F9F" => data <= "0000000000";
                when x"1FA0" => data <= "0000000000";
                when x"1FA1" => data <= "0000000000";
                when x"1FA2" => data <= "0000000000";
                when x"1FA3" => data <= "0000000000";
                when x"1FA4" => data <= "0000000000";
                when x"1FA5" => data <= "0000000000";
                when x"1FA6" => data <= "0000000000";
                when x"1FA7" => data <= "0000000000";
                when x"1FA8" => data <= "0000000000";
                when x"1FA9" => data <= "0000000000";
                when x"1FAA" => data <= "0000000000";
                when x"1FAB" => data <= "0000000000";
                when x"1FAC" => data <= "0000000000";
                when x"1FAD" => data <= "0000000000";
                when x"1FAE" => data <= "0000000000";
                when x"1FAF" => data <= "0000000000";
                when x"1FB0" => data <= "0000000000";
                when x"1FB1" => data <= "0000000000";
                when x"1FB2" => data <= "0000000000";
                when x"1FB3" => data <= "0000000000";
                when x"1FB4" => data <= "0000000000";
                when x"1FB5" => data <= "0000000000";
                when x"1FB6" => data <= "0000000000";
                when x"1FB7" => data <= "0000000000";
                when x"1FB8" => data <= "0000000000";
                when x"1FB9" => data <= "0000000000";
                when x"1FBA" => data <= "0000000000";
                when x"1FBB" => data <= "0000000000";
                when x"1FBC" => data <= "0000000000";
                when x"1FBD" => data <= "0000000000";
                when x"1FBE" => data <= "0000000000";
                when x"1FBF" => data <= "0000000000";
                when x"1FC0" => data <= "0000000000";
                when x"1FC1" => data <= "0000000000";
                when x"1FC2" => data <= "0000000000";
                when x"1FC3" => data <= "0000000000";
                when x"1FC4" => data <= "0000000000";
                when x"1FC5" => data <= "0000000000";
                when x"1FC6" => data <= "0000000000";
                when x"1FC7" => data <= "0000000000";
                when x"1FC8" => data <= "0000000000";
                when x"1FC9" => data <= "0000000000";
                when x"1FCA" => data <= "0000000000";
                when x"1FCB" => data <= "0000000000";
                when x"1FCC" => data <= "0000000000";
                when x"1FCD" => data <= "0000000000";
                when x"1FCE" => data <= "0000000000";
                when x"1FCF" => data <= "0000000000";
                when x"1FD0" => data <= "0000000000";
                when x"1FD1" => data <= "0000000000";
                when x"1FD2" => data <= "0000000000";
                when x"1FD3" => data <= "0000000000";
                when x"1FD4" => data <= "0000000000";
                when x"1FD5" => data <= "0000000000";
                when x"1FD6" => data <= "0000000000";
                when x"1FD7" => data <= "0000000000";
                when x"1FD8" => data <= "0000000000";
                when x"1FD9" => data <= "0000000000";
                when x"1FDA" => data <= "0000000000";
                when x"1FDB" => data <= "0000000000";
                when x"1FDC" => data <= "0000000000";
                when x"1FDD" => data <= "0000000000";
                when x"1FDE" => data <= "0000000000";
                when x"1FDF" => data <= "0000000000";
                when x"1FE0" => data <= "0000000000";
                when x"1FE1" => data <= "0000000000";
                when x"1FE2" => data <= "0000000000";
                when x"1FE3" => data <= "0000000000";
                when x"1FE4" => data <= "0000000000";
                when x"1FE5" => data <= "0000000000";
                when x"1FE6" => data <= "0000000000";
                when x"1FE7" => data <= "0000000000";
                when x"1FE8" => data <= "0000000000";
                when x"1FE9" => data <= "0000000000";
                when x"1FEA" => data <= "0000000000";
                when x"1FEB" => data <= "0000000000";
                when x"1FEC" => data <= "0000000000";
                when x"1FED" => data <= "0000000000";
                when x"1FEE" => data <= "0000000000";
                when x"1FEF" => data <= "0000000000";
                when x"1FF0" => data <= "0000000000";
                when x"1FF1" => data <= "0000000000";
                when x"1FF2" => data <= "0000000000";
                when x"1FF3" => data <= "0000000000";
                when x"1FF4" => data <= "0000000000";
                when x"1FF5" => data <= "0000000000";
                when x"1FF6" => data <= "0000000000";
                when x"1FF7" => data <= "0000000000";
                when x"1FF8" => data <= "0000000000";
                when x"1FF9" => data <= "0000000000";
                when x"1FFA" => data <= "0000000000";
                when x"1FFB" => data <= "0000000000";
                when x"1FFC" => data <= "0000000000";
                when x"1FFD" => data <= "0000000000";
                when x"1FFE" => data <= "0000000000";
                when x"1FFF" => data <= "0000000000";
                when x"2000" => data <= "0000000000";
                when x"2001" => data <= "0000000000";
                when x"2002" => data <= "0000000000";
                when x"2003" => data <= "0000000000";
                when x"2004" => data <= "0000000000";
                when x"2005" => data <= "0000000000";
                when x"2006" => data <= "0000000000";
                when x"2007" => data <= "0000000000";
                when x"2008" => data <= "0000000000";
                when x"2009" => data <= "0000000000";
                when x"200A" => data <= "0000000000";
                when x"200B" => data <= "0000000000";
                when x"200C" => data <= "0000000000";
                when x"200D" => data <= "0000000000";
                when x"200E" => data <= "0000000000";
                when x"200F" => data <= "0000000000";
                when x"2010" => data <= "0000000000";
                when x"2011" => data <= "0000000000";
                when x"2012" => data <= "0000000000";
                when x"2013" => data <= "0000000000";
                when x"2014" => data <= "0000000000";
                when x"2015" => data <= "0000000000";
                when x"2016" => data <= "0000000000";
                when x"2017" => data <= "0000000000";
                when x"2018" => data <= "0000000000";
                when x"2019" => data <= "0000000000";
                when x"201A" => data <= "0000000000";
                when x"201B" => data <= "0000000000";
                when x"201C" => data <= "0000000000";
                when x"201D" => data <= "0000000000";
                when x"201E" => data <= "0000000000";
                when x"201F" => data <= "0000000000";
                when x"2020" => data <= "0000000000";
                when x"2021" => data <= "0000000000";
                when x"2022" => data <= "0000000000";
                when x"2023" => data <= "0000000000";
                when x"2024" => data <= "1111011011";
                when x"2025" => data <= "0000000000";
                when x"2026" => data <= "0000000000";
                when x"2027" => data <= "0000000000";
                when x"2028" => data <= "0000000000";
                when x"2029" => data <= "0000000000";
                when x"202A" => data <= "0000000000";
                when x"202B" => data <= "0000000000";
                when x"202C" => data <= "0000000000";
                when x"202D" => data <= "0000000000";
                when x"202E" => data <= "0000000000";
                when x"202F" => data <= "0000000000";
                when x"2030" => data <= "0000000000";
                when x"2031" => data <= "0000000000";
                when x"2032" => data <= "0000000000";
                when x"2033" => data <= "0000000000";
                when x"2034" => data <= "0000000000";
                when x"2035" => data <= "0000000000";
                when x"2036" => data <= "0000000000";
                when x"2037" => data <= "0000000000";
                when x"2038" => data <= "0000000000";
                when x"2039" => data <= "0000000000";
                when x"203A" => data <= "0000000000";
                when x"203B" => data <= "0000000000";
                when x"203C" => data <= "0000000000";
                when x"203D" => data <= "0000000000";
                when x"203E" => data <= "0000000000";
                when x"203F" => data <= "0000000000";
                when x"2040" => data <= "0000000000";
                when x"2041" => data <= "0000000000";
                when x"2042" => data <= "0000000000";
                when x"2043" => data <= "0000000000";
                when x"2044" => data <= "0000000000";
                when x"2045" => data <= "0000000000";
                when x"2046" => data <= "0000000000";
                when x"2047" => data <= "0000000000";
                when x"2048" => data <= "0000000000";
                when x"2049" => data <= "0000000000";
                when x"204A" => data <= "0000000000";
                when x"204B" => data <= "0000000000";
                when x"204C" => data <= "0000000000";
                when x"204D" => data <= "0000000000";
                when x"204E" => data <= "0000000000";
                when x"204F" => data <= "0000000000";
                when x"2050" => data <= "0000000000";
                when x"2051" => data <= "0111110111";
                when x"2052" => data <= "0000000000";
                when x"2053" => data <= "0000000000";
                when x"2054" => data <= "0000000000";
                when x"2055" => data <= "0000000000";
                when x"2056" => data <= "0000000000";
                when x"2057" => data <= "0000000000";
                when x"2058" => data <= "0000000000";
                when x"2059" => data <= "0000000000";
                when x"205A" => data <= "0000000000";
                when x"205B" => data <= "0000000000";
                when x"205C" => data <= "0000000000";
                when x"205D" => data <= "0000000000";
                when x"205E" => data <= "0000000000";
                when x"205F" => data <= "0000000000";
                when x"2060" => data <= "0000000000";
                when x"2061" => data <= "0000000000";
                when x"2062" => data <= "0000000000";
                when x"2063" => data <= "0000000000";
                when x"2064" => data <= "0000000000";
                when x"2065" => data <= "0000000000";
                when x"2066" => data <= "0000000000";
                when x"2067" => data <= "0000000000";
                when x"2068" => data <= "0000000000";
                when x"2069" => data <= "0000000000";
                when x"206A" => data <= "0000000000";
                when x"206B" => data <= "0000000000";
                when x"206C" => data <= "0000000000";
                when x"206D" => data <= "0000000000";
                when x"206E" => data <= "0000000000";
                when x"206F" => data <= "0000000000";
                when x"2070" => data <= "0000000000";
                when x"2071" => data <= "0000000000";
                when x"2072" => data <= "0000000000";
                when x"2073" => data <= "0000000000";
                when x"2074" => data <= "0000000000";
                when x"2075" => data <= "0000000000";
                when x"2076" => data <= "0000000000";
                when x"2077" => data <= "0000000000";
                when x"2078" => data <= "0000000000";
                when x"2079" => data <= "0000000000";
                when x"207A" => data <= "0000000000";
                when x"207B" => data <= "0000000000";
                when x"207C" => data <= "0000000000";
                when x"207D" => data <= "0000000000";
                when x"207E" => data <= "0000000000";
                when x"207F" => data <= "0000000000";
                when x"2080" => data <= "0000000000";
                when x"2081" => data <= "0000000000";
                when x"2082" => data <= "0000000000";
                when x"2083" => data <= "0000000000";
                when x"2084" => data <= "0000000000";
                when x"2085" => data <= "0000000000";
                when x"2086" => data <= "0000000000";
                when x"2087" => data <= "0000000000";
                when x"2088" => data <= "0000000000";
                when x"2089" => data <= "0000000000";
                when x"208A" => data <= "0000000000";
                when x"208B" => data <= "0000000000";
                when x"208C" => data <= "0000000000";
                when x"208D" => data <= "0000000000";
                when x"208E" => data <= "0000000000";
                when x"208F" => data <= "0000000000";
                when x"2090" => data <= "0000000000";
                when x"2091" => data <= "0000000000";
                when x"2092" => data <= "0000000000";
                when x"2093" => data <= "0000000000";
                when x"2094" => data <= "0000000000";
                when x"2095" => data <= "0000000000";
                when x"2096" => data <= "0000000000";
                when x"2097" => data <= "0000000000";
                when x"2098" => data <= "0000000000";
                when x"2099" => data <= "0000000000";
                when x"209A" => data <= "0000000000";
                when x"209B" => data <= "0000000000";
                when x"209C" => data <= "0000000000";
                when x"209D" => data <= "0000000000";
                when x"209E" => data <= "0000000000";
                when x"209F" => data <= "0000000000";
                when x"20A0" => data <= "0000000000";
                when x"20A1" => data <= "0000000000";
                when x"20A2" => data <= "0000000000";
                when x"20A3" => data <= "0000000000";
                when x"20A4" => data <= "0000000000";
                when x"20A5" => data <= "0000000000";
                when x"20A6" => data <= "0000000000";
                when x"20A7" => data <= "0000000000";
                when x"20A8" => data <= "0000000000";
                when x"20A9" => data <= "0000000000";
                when x"20AA" => data <= "0000000000";
                when x"20AB" => data <= "0000000000";
                when x"20AC" => data <= "0000000000";
                when x"20AD" => data <= "0000000000";
                when x"20AE" => data <= "0000000000";
                when x"20AF" => data <= "0000000000";
                when x"20B0" => data <= "0000000000";
                when x"20B1" => data <= "0000000000";
                when x"20B2" => data <= "0000000000";
                when x"20B3" => data <= "0000000000";
                when x"20B4" => data <= "0000000000";
                when x"20B5" => data <= "0000000000";
                when x"20B6" => data <= "0000000000";
                when x"20B7" => data <= "0000000000";
                when x"20B8" => data <= "0000000000";
                when x"20B9" => data <= "0000000000";
                when x"20BA" => data <= "0000000000";
                when x"20BB" => data <= "0000000000";
                when x"20BC" => data <= "0000000000";
                when x"20BD" => data <= "0000000000";
                when x"20BE" => data <= "0000000000";
                when x"20BF" => data <= "0000000000";
                when x"20C0" => data <= "0000000000";
                when x"20C1" => data <= "0000000000";
                when x"20C2" => data <= "0000000000";
                when x"20C3" => data <= "0000000000";
                when x"20C4" => data <= "0000000000";
                when x"20C5" => data <= "0000000000";
                when x"20C6" => data <= "0000000000";
                when x"20C7" => data <= "0000000000";
                when x"20C8" => data <= "0000000000";
                when x"20C9" => data <= "0000000000";
                when x"20CA" => data <= "0000000000";
                when x"20CB" => data <= "0000000000";
                when x"20CC" => data <= "0000000000";
                when x"20CD" => data <= "0000000000";
                when x"20CE" => data <= "0000000000";
                when x"20CF" => data <= "0000000000";
                when x"20D0" => data <= "0000000000";
                when x"20D1" => data <= "0000000000";
                when x"20D2" => data <= "0000000000";
                when x"20D3" => data <= "0000000000";
                when x"20D4" => data <= "0000000000";
                when x"20D5" => data <= "0000000000";
                when x"20D6" => data <= "0000000000";
                when x"20D7" => data <= "0000000000";
                when x"20D8" => data <= "0000000000";
                when x"20D9" => data <= "0000000000";
                when x"20DA" => data <= "0000000000";
                when x"20DB" => data <= "0000000000";
                when x"20DC" => data <= "0000000000";
                when x"20DD" => data <= "0000000000";
                when x"20DE" => data <= "0000000000";
                when x"20DF" => data <= "0000000000";
                when x"20E0" => data <= "0000000000";
                when x"20E1" => data <= "0000000000";
                when x"20E2" => data <= "0000000000";
                when x"20E3" => data <= "0000000000";
                when x"20E4" => data <= "0000000000";
                when x"20E5" => data <= "0000000000";
                when x"20E6" => data <= "0000000000";
                when x"20E7" => data <= "0000000000";
                when x"20E8" => data <= "0000000000";
                when x"20E9" => data <= "0000000000";
                when x"20EA" => data <= "0000000000";
                when x"20EB" => data <= "0000000000";
                when x"20EC" => data <= "0000000000";
                when x"20ED" => data <= "0000000000";
                when x"20EE" => data <= "0000000000";
                when x"20EF" => data <= "0000000000";
                when x"20F0" => data <= "0000000000";
                when x"20F1" => data <= "0000000000";
                when x"20F2" => data <= "0000000000";
                when x"20F3" => data <= "0000000000";
                when x"20F4" => data <= "0000000000";
                when x"20F5" => data <= "0000000000";
                when x"20F6" => data <= "0000000000";
                when x"20F7" => data <= "0000000000";
                when x"20F8" => data <= "0000000000";
                when x"20F9" => data <= "0000000000";
                when x"20FA" => data <= "0000000000";
                when x"20FB" => data <= "0000000000";
                when x"20FC" => data <= "0000000000";
                when x"20FD" => data <= "0000000000";
                when x"20FE" => data <= "0000000000";
                when x"20FF" => data <= "0000000000";
                when x"2100" => data <= "0000000000";
                when x"2101" => data <= "0000000000";
                when x"2102" => data <= "0000000000";
                when x"2103" => data <= "0000000000";
                when x"2104" => data <= "0000000000";
                when x"2105" => data <= "0000000000";
                when x"2106" => data <= "0000000000";
                when x"2107" => data <= "0000000000";
                when x"2108" => data <= "0000000000";
                when x"2109" => data <= "0000000000";
                when x"210A" => data <= "0000000000";
                when x"210B" => data <= "0000000000";
                when x"210C" => data <= "0000000000";
                when x"210D" => data <= "0000000000";
                when x"210E" => data <= "0000000000";
                when x"210F" => data <= "0000000000";
                when x"2110" => data <= "0000000000";
                when x"2111" => data <= "0000000000";
                when x"2112" => data <= "0000000000";
                when x"2113" => data <= "0000000000";
                when x"2114" => data <= "0000000000";
                when x"2115" => data <= "0000000000";
                when x"2116" => data <= "0000000000";
                when x"2117" => data <= "0000000000";
                when x"2118" => data <= "0000000000";
                when x"2119" => data <= "0000000000";
                when x"211A" => data <= "0000000000";
                when x"211B" => data <= "0000000000";
                when x"211C" => data <= "0000000000";
                when x"211D" => data <= "0000000000";
                when x"211E" => data <= "0000000000";
                when x"211F" => data <= "0000000000";
                when x"2120" => data <= "0000000000";
                when x"2121" => data <= "0000000000";
                when x"2122" => data <= "0000000000";
                when x"2123" => data <= "0000000000";
                when x"2124" => data <= "0000000000";
                when x"2125" => data <= "0000000000";
                when x"2126" => data <= "0000000000";
                when x"2127" => data <= "0000000000";
                when x"2128" => data <= "0000000000";
                when x"2129" => data <= "0000000000";
                when x"212A" => data <= "0000000000";
                when x"212B" => data <= "0000000000";
                when x"212C" => data <= "0000000000";
                when x"212D" => data <= "0000000000";
                when x"212E" => data <= "0000000000";
                when x"212F" => data <= "0000000000";
                when x"2130" => data <= "0000000000";
                when x"2131" => data <= "0000000000";
                when x"2132" => data <= "0000000000";
                when x"2133" => data <= "0000000000";
                when x"2134" => data <= "0000000000";
                when x"2135" => data <= "0000000000";
                when x"2136" => data <= "0000000000";
                when x"2137" => data <= "0000000000";
                when x"2138" => data <= "0000000000";
                when x"2139" => data <= "0000000000";
                when x"213A" => data <= "0000000000";
                when x"213B" => data <= "0000000000";
                when x"213C" => data <= "0000000000";
                when x"213D" => data <= "0000000000";
                when x"213E" => data <= "0000000000";
                when x"213F" => data <= "0000000000";
                when x"2140" => data <= "0000000000";
                when x"2141" => data <= "0000000000";
                when x"2142" => data <= "0000000000";
                when x"2143" => data <= "0000000000";
                when x"2144" => data <= "0000000000";
                when x"2145" => data <= "0000000000";
                when x"2146" => data <= "0000000000";
                when x"2147" => data <= "0000000000";
                when x"2148" => data <= "0000000000";
                when x"2149" => data <= "0000000000";
                when x"214A" => data <= "0000000000";
                when x"214B" => data <= "0000000000";
                when x"214C" => data <= "0000000000";
                when x"214D" => data <= "0000000000";
                when x"214E" => data <= "0000000000";
                when x"214F" => data <= "0000000000";
                when x"2150" => data <= "0000000000";
                when x"2151" => data <= "0000000000";
                when x"2152" => data <= "0000000000";
                when x"2153" => data <= "0000000000";
                when x"2154" => data <= "0000000000";
                when x"2155" => data <= "0000000000";
                when x"2156" => data <= "0000000000";
                when x"2157" => data <= "0000000000";
                when x"2158" => data <= "0000000000";
                when x"2159" => data <= "0000000000";
                when x"215A" => data <= "0000000000";
                when x"215B" => data <= "0000000000";
                when x"215C" => data <= "0000000000";
                when x"215D" => data <= "0000000000";
                when x"215E" => data <= "0000000000";
                when x"215F" => data <= "0000000000";
                when x"2160" => data <= "0000000000";
                when x"2161" => data <= "0000000000";
                when x"2162" => data <= "0000000000";
                when x"2163" => data <= "0000000000";
                when x"2164" => data <= "0000000000";
                when x"2165" => data <= "0000000000";
                when x"2166" => data <= "0000000000";
                when x"2167" => data <= "0000000000";
                when x"2168" => data <= "0000000000";
                when x"2169" => data <= "0000000000";
                when x"216A" => data <= "0000000000";
                when x"216B" => data <= "0000000000";
                when x"216C" => data <= "0000000000";
                when x"216D" => data <= "0000000000";
                when x"216E" => data <= "0000000000";
                when x"216F" => data <= "0000000000";
                when x"2170" => data <= "0000000000";
                when x"2171" => data <= "0000000000";
                when x"2172" => data <= "0000000000";
                when x"2173" => data <= "0000000000";
                when x"2174" => data <= "0000000000";
                when x"2175" => data <= "0000000000";
                when x"2176" => data <= "0000000000";
                when x"2177" => data <= "0000000000";
                when x"2178" => data <= "0000000000";
                when x"2179" => data <= "0000000000";
                when x"217A" => data <= "0000000000";
                when x"217B" => data <= "0000000000";
                when x"217C" => data <= "0000000000";
                when x"217D" => data <= "0000000000";
                when x"217E" => data <= "0000000000";
                when x"217F" => data <= "0000000000";
                when x"2180" => data <= "0000000000";
                when x"2181" => data <= "0000000000";
                when x"2182" => data <= "0000000000";
                when x"2183" => data <= "0000000000";
                when x"2184" => data <= "0000000000";
                when x"2185" => data <= "0000000000";
                when x"2186" => data <= "0111110111";
                when x"2187" => data <= "0000000000";
                when x"2188" => data <= "0000000000";
                when x"2189" => data <= "0000000000";
                when x"218A" => data <= "0000000000";
                when x"218B" => data <= "0000000000";
                when x"218C" => data <= "0000000000";
                when x"218D" => data <= "0000000000";
                when x"218E" => data <= "0000000000";
                when x"218F" => data <= "0000000000";
                when x"2190" => data <= "0000000000";
                when x"2191" => data <= "0000000000";
                when x"2192" => data <= "0000000000";
                when x"2193" => data <= "0000000000";
                when x"2194" => data <= "0000000000";
                when x"2195" => data <= "0000000000";
                when x"2196" => data <= "0000000000";
                when x"2197" => data <= "0000000000";
                when x"2198" => data <= "0000000000";
                when x"2199" => data <= "0000000000";
                when x"219A" => data <= "0000000000";
                when x"219B" => data <= "0000000000";
                when x"219C" => data <= "0000000000";
                when x"219D" => data <= "0000000000";
                when x"219E" => data <= "0000000000";
                when x"219F" => data <= "0000000000";
                when x"21A0" => data <= "0000000000";
                when x"21A1" => data <= "0000000000";
                when x"21A2" => data <= "0000000000";
                when x"21A3" => data <= "0000000000";
                when x"21A4" => data <= "0000000000";
                when x"21A5" => data <= "0000000000";
                when x"21A6" => data <= "0000000000";
                when x"21A7" => data <= "0000000000";
                when x"21A8" => data <= "0000000000";
                when x"21A9" => data <= "0000000000";
                when x"21AA" => data <= "0000000000";
                when x"21AB" => data <= "0000000000";
                when x"21AC" => data <= "0000000000";
                when x"21AD" => data <= "0000000000";
                when x"21AE" => data <= "0000000000";
                when x"21AF" => data <= "0000000000";
                when x"21B0" => data <= "0000000000";
                when x"21B1" => data <= "0000000000";
                when x"21B2" => data <= "0000000000";
                when x"21B3" => data <= "0000000000";
                when x"21B4" => data <= "0000000000";
                when x"21B5" => data <= "0000000000";
                when x"21B6" => data <= "0000000000";
                when x"21B7" => data <= "0000000000";
                when x"21B8" => data <= "0000000000";
                when x"21B9" => data <= "0000000000";
                when x"21BA" => data <= "0000000000";
                when x"21BB" => data <= "0000000000";
                when x"21BC" => data <= "0000000000";
                when x"21BD" => data <= "0000000000";
                when x"21BE" => data <= "0000000000";
                when x"21BF" => data <= "0000000000";
                when x"21C0" => data <= "0000000000";
                when x"21C1" => data <= "0000000000";
                when x"21C2" => data <= "0000000000";
                when x"21C3" => data <= "0000000000";
                when x"21C4" => data <= "0000000000";
                when x"21C5" => data <= "0000000000";
                when x"21C6" => data <= "0000000000";
                when x"21C7" => data <= "0000000000";
                when x"21C8" => data <= "0000000000";
                when x"21C9" => data <= "0000000000";
                when x"21CA" => data <= "0000000000";
                when x"21CB" => data <= "0000000000";
                when x"21CC" => data <= "0000000000";
                when x"21CD" => data <= "0000000000";
                when x"21CE" => data <= "0000000000";
                when x"21CF" => data <= "0000000000";
                when x"21D0" => data <= "0000000000";
                when x"21D1" => data <= "0000000000";
                when x"21D2" => data <= "0000000000";
                when x"21D3" => data <= "0000000000";
                when x"21D4" => data <= "0000000000";
                when x"21D5" => data <= "0000000000";
                when x"21D6" => data <= "0000000000";
                when x"21D7" => data <= "0000000000";
                when x"21D8" => data <= "0000000000";
                when x"21D9" => data <= "0000000000";
                when x"21DA" => data <= "0000000000";
                when x"21DB" => data <= "0000000000";
                when x"21DC" => data <= "0000000000";
                when x"21DD" => data <= "0000000000";
                when x"21DE" => data <= "0000000000";
                when x"21DF" => data <= "0000000000";
                when x"21E0" => data <= "0000000000";
                when x"21E1" => data <= "0000000000";
                when x"21E2" => data <= "0000000000";
                when x"21E3" => data <= "0000000000";
                when x"21E4" => data <= "0000000000";
                when x"21E5" => data <= "0000000000";
                when x"21E6" => data <= "1111011011";
                when x"21E7" => data <= "0000000000";
                when x"21E8" => data <= "0000000000";
                when x"21E9" => data <= "0000000000";
                when x"21EA" => data <= "0000000000";
                when x"21EB" => data <= "0000000000";
                when x"21EC" => data <= "0000000000";
                when x"21ED" => data <= "0000000000";
                when x"21EE" => data <= "0000000000";
                when x"21EF" => data <= "0000000000";
                when x"21F0" => data <= "0000000000";
                when x"21F1" => data <= "0000000000";
                when x"21F2" => data <= "0000000000";
                when x"21F3" => data <= "0000000000";
                when x"21F4" => data <= "0000000000";
                when x"21F5" => data <= "0000000000";
                when x"21F6" => data <= "0000000000";
                when x"21F7" => data <= "0000000000";
                when x"21F8" => data <= "0000000000";
                when x"21F9" => data <= "0000000000";
                when x"21FA" => data <= "0000000000";
                when x"21FB" => data <= "0000000000";
                when x"21FC" => data <= "0000000000";
                when x"21FD" => data <= "0000000000";
                when x"21FE" => data <= "0000000000";
                when x"21FF" => data <= "0000000000";
                when x"2200" => data <= "0000000000";
                when x"2201" => data <= "0000000000";
                when x"2202" => data <= "0000000000";
                when x"2203" => data <= "0000000000";
                when x"2204" => data <= "0000000000";
                when x"2205" => data <= "0000000000";
                when x"2206" => data <= "0000000000";
                when x"2207" => data <= "0000000000";
                when x"2208" => data <= "0000000000";
                when x"2209" => data <= "0000000000";
                when x"220A" => data <= "0000000000";
                when x"220B" => data <= "0000000000";
                when x"220C" => data <= "0000000000";
                when x"220D" => data <= "0000000000";
                when x"220E" => data <= "0000000000";
                when x"220F" => data <= "0000000000";
                when x"2210" => data <= "0000000000";
                when x"2211" => data <= "0000000000";
                when x"2212" => data <= "0000000000";
                when x"2213" => data <= "0000000000";
                when x"2214" => data <= "0000000000";
                when x"2215" => data <= "0000000000";
                when x"2216" => data <= "0000000000";
                when x"2217" => data <= "0000000000";
                when x"2218" => data <= "0000000000";
                when x"2219" => data <= "0000000000";
                when x"221A" => data <= "0000000000";
                when x"221B" => data <= "0000000000";
                when x"221C" => data <= "0000000000";
                when x"221D" => data <= "0000000000";
                when x"221E" => data <= "0000000000";
                when x"221F" => data <= "0000000000";
                when x"2220" => data <= "0111110111";
                when x"2221" => data <= "0000000000";
                when x"2222" => data <= "0000000000";
                when x"2223" => data <= "0111110111";
                when x"2224" => data <= "0000000000";
                when x"2225" => data <= "0000000000";
                when x"2226" => data <= "0000000000";
                when x"2227" => data <= "0000000000";
                when x"2228" => data <= "1101010000";
                when x"2229" => data <= "0000000000";
                when x"222A" => data <= "0000000000";
                when x"222B" => data <= "0000000000";
                when x"222C" => data <= "0000000000";
                when x"222D" => data <= "0000000000";
                when x"222E" => data <= "0000000000";
                when x"222F" => data <= "0000000000";
                when x"2230" => data <= "0000000000";
                when x"2231" => data <= "0000000000";
                when x"2232" => data <= "0000000000";
                when x"2233" => data <= "0000000000";
                when x"2234" => data <= "0000000000";
                when x"2235" => data <= "0000000000";
                when x"2236" => data <= "0000000000";
                when x"2237" => data <= "0000000000";
                when x"2238" => data <= "0000000000";
                when x"2239" => data <= "0000000000";
                when x"223A" => data <= "0000000000";
                when x"223B" => data <= "0000000000";
                when x"223C" => data <= "0000000000";
                when x"223D" => data <= "0000000000";
                when x"223E" => data <= "0000000000";
                when x"223F" => data <= "0000000000";
                when x"2240" => data <= "0000000000";
                when x"2241" => data <= "0000000000";
                when x"2242" => data <= "0000000000";
                when x"2243" => data <= "0000000000";
                when x"2244" => data <= "0000000000";
                when x"2245" => data <= "0000000000";
                when x"2246" => data <= "0000000000";
                when x"2247" => data <= "0000000000";
                when x"2248" => data <= "0000000000";
                when x"2249" => data <= "0000000000";
                when x"224A" => data <= "0000000000";
                when x"224B" => data <= "0000000000";
                when x"224C" => data <= "0000000000";
                when x"224D" => data <= "0000000000";
                when x"224E" => data <= "0000000000";
                when x"224F" => data <= "0000000000";
                when x"2250" => data <= "0000000000";
                when x"2251" => data <= "0000000000";
                when x"2252" => data <= "0000000000";
                when x"2253" => data <= "0000000000";
                when x"2254" => data <= "0000000000";
                when x"2255" => data <= "0000000000";
                when x"2256" => data <= "0000000000";
                when x"2257" => data <= "0000000000";
                when x"2258" => data <= "0000000000";
                when x"2259" => data <= "0000000000";
                when x"225A" => data <= "0000000000";
                when x"225B" => data <= "0000000000";
                when x"225C" => data <= "0000000000";
                when x"225D" => data <= "0000000000";
                when x"225E" => data <= "0000000000";
                when x"225F" => data <= "0000000000";
                when x"2260" => data <= "0000000000";
                when x"2261" => data <= "0000000000";
                when x"2262" => data <= "0000000000";
                when x"2263" => data <= "0000000000";
                when x"2264" => data <= "0000000000";
                when x"2265" => data <= "0000000000";
                when x"2266" => data <= "0000000000";
                when x"2267" => data <= "0000000000";
                when x"2268" => data <= "1101010000";
                when x"2269" => data <= "0000000000";
                when x"226A" => data <= "0000000000";
                when x"226B" => data <= "0000000000";
                when x"226C" => data <= "0000000000";
                when x"226D" => data <= "0000000000";
                when x"226E" => data <= "0000000000";
                when x"226F" => data <= "0000000000";
                when x"2270" => data <= "0000000000";
                when x"2271" => data <= "0000000000";
                when x"2272" => data <= "0000000000";
                when x"2273" => data <= "0000000000";
                when x"2274" => data <= "0000000000";
                when x"2275" => data <= "0000000000";
                when x"2276" => data <= "0000000000";
                when x"2277" => data <= "0000000000";
                when x"2278" => data <= "0000000000";
                when x"2279" => data <= "0000000000";
                when x"227A" => data <= "0000000000";
                when x"227B" => data <= "0000000000";
                when x"227C" => data <= "0000000000";
                when x"227D" => data <= "0000000000";
                when x"227E" => data <= "0000000000";
                when x"227F" => data <= "0000000000";
                when x"2280" => data <= "0000000000";
                when x"2281" => data <= "0000000000";
                when x"2282" => data <= "0000000000";
                when x"2283" => data <= "0000000000";
                when x"2284" => data <= "0000000000";
                when x"2285" => data <= "0000000000";
                when x"2286" => data <= "0000000000";
                when x"2287" => data <= "0000000000";
                when x"2288" => data <= "0000000000";
                when x"2289" => data <= "0000000000";
                when x"228A" => data <= "0000000000";
                when x"228B" => data <= "0000000000";
                when x"228C" => data <= "0000000000";
                when x"228D" => data <= "0000000000";
                when x"228E" => data <= "0000000000";
                when x"228F" => data <= "0000000000";
                when x"2290" => data <= "0000000000";
                when x"2291" => data <= "0000000000";
                when x"2292" => data <= "0000000000";
                when x"2293" => data <= "0000000000";
                when x"2294" => data <= "0000000000";
                when x"2295" => data <= "0000000000";
                when x"2296" => data <= "0000000000";
                when x"2297" => data <= "0000000000";
                when x"2298" => data <= "0000000000";
                when x"2299" => data <= "0000000000";
                when x"229A" => data <= "0000000000";
                when x"229B" => data <= "0000000000";
                when x"229C" => data <= "0000000000";
                when x"229D" => data <= "0000000000";
                when x"229E" => data <= "0000000000";
                when x"229F" => data <= "0000000000";
                when x"22A0" => data <= "0000000000";
                when x"22A1" => data <= "0000000000";
                when x"22A2" => data <= "0000000000";
                when x"22A3" => data <= "0000000000";
                when x"22A4" => data <= "0000000000";
                when x"22A5" => data <= "0000000000";
                when x"22A6" => data <= "0000000000";
                when x"22A7" => data <= "0000000000";
                when x"22A8" => data <= "0000000000";
                when x"22A9" => data <= "0000000000";
                when x"22AA" => data <= "0000000000";
                when x"22AB" => data <= "0000000000";
                when x"22AC" => data <= "0000000000";
                when x"22AD" => data <= "0000000000";
                when x"22AE" => data <= "0000000000";
                when x"22AF" => data <= "0000000000";
                when x"22B0" => data <= "0000000000";
                when x"22B1" => data <= "0000000000";
                when x"22B2" => data <= "0000000000";
                when x"22B3" => data <= "0000000000";
                when x"22B4" => data <= "0000000000";
                when x"22B5" => data <= "0000000000";
                when x"22B6" => data <= "0000000000";
                when x"22B7" => data <= "0000000000";
                when x"22B8" => data <= "0000000000";
                when x"22B9" => data <= "0000000000";
                when x"22BA" => data <= "0000000000";
                when x"22BB" => data <= "0000000000";
                when x"22BC" => data <= "0000000000";
                when x"22BD" => data <= "0000000000";
                when x"22BE" => data <= "0000000000";
                when x"22BF" => data <= "0000000000";
                when x"22C0" => data <= "0000000000";
                when x"22C1" => data <= "0000000000";
                when x"22C2" => data <= "0000000000";
                when x"22C3" => data <= "0000000000";
                when x"22C4" => data <= "0000000000";
                when x"22C5" => data <= "0000000000";
                when x"22C6" => data <= "0000000000";
                when x"22C7" => data <= "0000000000";
                when x"22C8" => data <= "0000000000";
                when x"22C9" => data <= "0000000000";
                when x"22CA" => data <= "0000000000";
                when x"22CB" => data <= "0000000000";
                when x"22CC" => data <= "0000000000";
                when x"22CD" => data <= "0000000000";
                when x"22CE" => data <= "0000000000";
                when x"22CF" => data <= "0000000000";
                when x"22D0" => data <= "0000000000";
                when x"22D1" => data <= "0000000000";
                when x"22D2" => data <= "0000000000";
                when x"22D3" => data <= "0000000000";
                when x"22D4" => data <= "0000000000";
                when x"22D5" => data <= "0000000000";
                when x"22D6" => data <= "0000000000";
                when x"22D7" => data <= "0000000000";
                when x"22D8" => data <= "0000000000";
                when x"22D9" => data <= "0000000000";
                when x"22DA" => data <= "0000000000";
                when x"22DB" => data <= "0000000000";
                when x"22DC" => data <= "0000000000";
                when x"22DD" => data <= "0000000000";
                when x"22DE" => data <= "0000000000";
                when x"22DF" => data <= "0000000000";
                when x"22E0" => data <= "0000000000";
                when x"22E1" => data <= "0000000000";
                when x"22E2" => data <= "0000000000";
                when x"22E3" => data <= "0000000000";
                when x"22E4" => data <= "0000000000";
                when x"22E5" => data <= "0000000000";
                when x"22E6" => data <= "0000000000";
                when x"22E7" => data <= "0000000000";
                when x"22E8" => data <= "0000000000";
                when x"22E9" => data <= "0000000000";
                when x"22EA" => data <= "0000000000";
                when x"22EB" => data <= "0000000000";
                when x"22EC" => data <= "0000000000";
                when x"22ED" => data <= "0000000000";
                when x"22EE" => data <= "0000000000";
                when x"22EF" => data <= "0000000000";
                when x"22F0" => data <= "0000000000";
                when x"22F1" => data <= "0000000000";
                when x"22F2" => data <= "0000000000";
                when x"22F3" => data <= "0000000000";
                when x"22F4" => data <= "0000000000";
                when x"22F5" => data <= "0000000000";
                when x"22F6" => data <= "0000000000";
                when x"22F7" => data <= "0000000000";
                when x"22F8" => data <= "0000000000";
                when x"22F9" => data <= "0000000000";
                when x"22FA" => data <= "0000000000";
                when x"22FB" => data <= "0000000000";
                when x"22FC" => data <= "0000000000";
                when x"22FD" => data <= "0000000000";
                when x"22FE" => data <= "0000000000";
                when x"22FF" => data <= "0000000000";
                when x"2300" => data <= "0000000000";
                when x"2301" => data <= "0000000000";
                when x"2302" => data <= "0000000000";
                when x"2303" => data <= "0000000000";
                when x"2304" => data <= "0000000000";
                when x"2305" => data <= "0000000000";
                when x"2306" => data <= "0000000000";
                when x"2307" => data <= "0000000000";
                when x"2308" => data <= "0000000000";
                when x"2309" => data <= "0000000000";
                when x"230A" => data <= "0000000000";
                when x"230B" => data <= "0000000000";
                when x"230C" => data <= "0000000000";
                when x"230D" => data <= "0000000000";
                when x"230E" => data <= "0000000000";
                when x"230F" => data <= "0000000000";
                when x"2310" => data <= "0000000000";
                when x"2311" => data <= "0000000000";
                when x"2312" => data <= "0000000000";
                when x"2313" => data <= "0000000000";
                when x"2314" => data <= "0000000000";
                when x"2315" => data <= "0000000000";
                when x"2316" => data <= "0000000000";
                when x"2317" => data <= "0000000000";
                when x"2318" => data <= "0000000000";
                when x"2319" => data <= "0000000000";
                when x"231A" => data <= "0000000000";
                when x"231B" => data <= "0000000000";
                when x"231C" => data <= "0000000000";
                when x"231D" => data <= "0000000000";
                when x"231E" => data <= "0000000000";
                when x"231F" => data <= "0000000000";
                when x"2320" => data <= "0000000000";
                when x"2321" => data <= "0000000000";
                when x"2322" => data <= "0000000000";
                when x"2323" => data <= "0000000000";
                when x"2324" => data <= "0000000000";
                when x"2325" => data <= "0000000000";
                when x"2326" => data <= "0000000000";
                when x"2327" => data <= "0000000000";
                when x"2328" => data <= "0000000000";
                when x"2329" => data <= "0000000000";
                when x"232A" => data <= "0000000000";
                when x"232B" => data <= "0000000000";
                when x"232C" => data <= "0000000000";
                when x"232D" => data <= "0000000000";
                when x"232E" => data <= "0000000000";
                when x"232F" => data <= "0000000000";
                when x"2330" => data <= "0000000000";
                when x"2331" => data <= "0000000000";
                when x"2332" => data <= "0000000000";
                when x"2333" => data <= "0000000000";
                when x"2334" => data <= "0000000000";
                when x"2335" => data <= "0000000000";
                when x"2336" => data <= "0000000000";
                when x"2337" => data <= "0000000000";
                when x"2338" => data <= "0000000000";
                when x"2339" => data <= "0000000000";
                when x"233A" => data <= "0000000000";
                when x"233B" => data <= "0000000000";
                when x"233C" => data <= "0000000000";
                when x"233D" => data <= "0000000000";
                when x"233E" => data <= "0000000000";
                when x"233F" => data <= "0000000000";
                when x"2340" => data <= "0000000000";
                when x"2341" => data <= "0000000000";
                when x"2342" => data <= "0000000000";
                when x"2343" => data <= "0000000000";
                when x"2344" => data <= "0000000000";
                when x"2345" => data <= "0000000000";
                when x"2346" => data <= "0000000000";
                when x"2347" => data <= "0000000000";
                when x"2348" => data <= "0000000000";
                when x"2349" => data <= "0000000000";
                when x"234A" => data <= "0000000000";
                when x"234B" => data <= "0000000000";
                when x"234C" => data <= "0000000000";
                when x"234D" => data <= "0000000000";
                when x"234E" => data <= "0000000000";
                when x"234F" => data <= "0000000000";
                when x"2350" => data <= "0000000000";
                when x"2351" => data <= "0000000000";
                when x"2352" => data <= "0000000000";
                when x"2353" => data <= "0000000000";
                when x"2354" => data <= "0000000000";
                when x"2355" => data <= "0000000000";
                when x"2356" => data <= "0000000000";
                when x"2357" => data <= "0111110111";
                when x"2358" => data <= "0000000000";
                when x"2359" => data <= "0000000000";
                when x"235A" => data <= "0000000000";
                when x"235B" => data <= "0000000000";
                when x"235C" => data <= "0000000000";
                when x"235D" => data <= "0000000000";
                when x"235E" => data <= "0000000000";
                when x"235F" => data <= "0000000000";
                when x"2360" => data <= "0000000000";
                when x"2361" => data <= "0000000000";
                when x"2362" => data <= "0000000000";
                when x"2363" => data <= "0000000000";
                when x"2364" => data <= "0000000000";
                when x"2365" => data <= "0000000000";
                when x"2366" => data <= "0000000000";
                when x"2367" => data <= "0000000000";
                when x"2368" => data <= "0000000000";
                when x"2369" => data <= "0000000000";
                when x"236A" => data <= "0000000000";
                when x"236B" => data <= "0000000000";
                when x"236C" => data <= "0000000000";
                when x"236D" => data <= "0000000000";
                when x"236E" => data <= "0000000000";
                when x"236F" => data <= "0000000000";
                when x"2370" => data <= "0000000000";
                when x"2371" => data <= "0000000000";
                when x"2372" => data <= "0000000000";
                when x"2373" => data <= "0000000000";
                when x"2374" => data <= "0000000000";
                when x"2375" => data <= "0000000000";
                when x"2376" => data <= "0000000000";
                when x"2377" => data <= "0000000000";
                when x"2378" => data <= "0000000000";
                when x"2379" => data <= "0000000000";
                when x"237A" => data <= "0000000000";
                when x"237B" => data <= "0000000000";
                when x"237C" => data <= "0000000000";
                when x"237D" => data <= "0000000000";
                when x"237E" => data <= "0000000000";
                when x"237F" => data <= "0000000000";
                when x"2380" => data <= "0000000000";
                when x"2381" => data <= "0000000000";
                when x"2382" => data <= "0000000000";
                when x"2383" => data <= "0000000000";
                when x"2384" => data <= "0000000000";
                when x"2385" => data <= "1100111010";
                when x"2386" => data <= "0000000000";
                when x"2387" => data <= "0000000000";
                when x"2388" => data <= "0000000000";
                when x"2389" => data <= "0000000000";
                when x"238A" => data <= "0000000000";
                when x"238B" => data <= "0000000000";
                when x"238C" => data <= "0000000000";
                when x"238D" => data <= "0000000000";
                when x"238E" => data <= "0000000000";
                when x"238F" => data <= "0000000000";
                when x"2390" => data <= "0000000000";
                when x"2391" => data <= "0000000000";
                when x"2392" => data <= "0000000000";
                when x"2393" => data <= "0000000000";
                when x"2394" => data <= "0000000000";
                when x"2395" => data <= "0000000000";
                when x"2396" => data <= "0000000000";
                when x"2397" => data <= "0000000000";
                when x"2398" => data <= "0000000000";
                when x"2399" => data <= "0000000000";
                when x"239A" => data <= "0000000000";
                when x"239B" => data <= "0000000000";
                when x"239C" => data <= "0000000000";
                when x"239D" => data <= "0000000000";
                when x"239E" => data <= "0000000000";
                when x"239F" => data <= "0000000000";
                when x"23A0" => data <= "0000000000";
                when x"23A1" => data <= "0000000000";
                when x"23A2" => data <= "0000000000";
                when x"23A3" => data <= "0000000000";
                when x"23A4" => data <= "0000000000";
                when x"23A5" => data <= "0000000000";
                when x"23A6" => data <= "0000000000";
                when x"23A7" => data <= "0000000000";
                when x"23A8" => data <= "0000000000";
                when x"23A9" => data <= "0000000000";
                when x"23AA" => data <= "0000000000";
                when x"23AB" => data <= "0000000000";
                when x"23AC" => data <= "0000000000";
                when x"23AD" => data <= "0000000000";
                when x"23AE" => data <= "0000000000";
                when x"23AF" => data <= "0000000000";
                when x"23B0" => data <= "0000000000";
                when x"23B1" => data <= "0000000000";
                when x"23B2" => data <= "0000000000";
                when x"23B3" => data <= "0000000000";
                when x"23B4" => data <= "0000000000";
                when x"23B5" => data <= "0000000000";
                when x"23B6" => data <= "0000000000";
                when x"23B7" => data <= "0000000000";
                when x"23B8" => data <= "0000000000";
                when x"23B9" => data <= "0000000000";
                when x"23BA" => data <= "0000000000";
                when x"23BB" => data <= "0000000000";
                when x"23BC" => data <= "0000000000";
                when x"23BD" => data <= "0000000000";
                when x"23BE" => data <= "0000000000";
                when x"23BF" => data <= "0000000000";
                when x"23C0" => data <= "0000000000";
                when x"23C1" => data <= "0000000000";
                when x"23C2" => data <= "0000000000";
                when x"23C3" => data <= "0000000000";
                when x"23C4" => data <= "0000000000";
                when x"23C5" => data <= "0000000000";
                when x"23C6" => data <= "0000000000";
                when x"23C7" => data <= "0000000000";
                when x"23C8" => data <= "0000000000";
                when x"23C9" => data <= "0000000000";
                when x"23CA" => data <= "0000000000";
                when x"23CB" => data <= "0000000000";
                when x"23CC" => data <= "0000000000";
                when x"23CD" => data <= "0000000000";
                when x"23CE" => data <= "0000000000";
                when x"23CF" => data <= "0000000000";
                when x"23D0" => data <= "0000000000";
                when x"23D1" => data <= "0000000000";
                when x"23D2" => data <= "0000000000";
                when x"23D3" => data <= "0000000000";
                when x"23D4" => data <= "0000000000";
                when x"23D5" => data <= "0000000000";
                when x"23D6" => data <= "0000000000";
                when x"23D7" => data <= "0000000000";
                when x"23D8" => data <= "0000000000";
                when x"23D9" => data <= "0000000000";
                when x"23DA" => data <= "0000000000";
                when x"23DB" => data <= "0000000000";
                when x"23DC" => data <= "0000000000";
                when x"23DD" => data <= "0000000000";
                when x"23DE" => data <= "0000000000";
                when x"23DF" => data <= "0000000000";
                when x"23E0" => data <= "0000000000";
                when x"23E1" => data <= "0000000000";
                when x"23E2" => data <= "0000000000";
                when x"23E3" => data <= "0000000000";
                when x"23E4" => data <= "0000000000";
                when x"23E5" => data <= "0000000000";
                when x"23E6" => data <= "0000000000";
                when x"23E7" => data <= "0000000000";
                when x"23E8" => data <= "0000000000";
                when x"23E9" => data <= "0000000000";
                when x"23EA" => data <= "0000000000";
                when x"23EB" => data <= "0000000000";
                when x"23EC" => data <= "0000000000";
                when x"23ED" => data <= "0000000000";
                when x"23EE" => data <= "0000000000";
                when x"23EF" => data <= "0000000000";
                when x"23F0" => data <= "0000000000";
                when x"23F1" => data <= "0000000000";
                when x"23F2" => data <= "0000000000";
                when x"23F3" => data <= "0000000000";
                when x"23F4" => data <= "0000000000";
                when x"23F5" => data <= "0000000000";
                when x"23F6" => data <= "0000000000";
                when x"23F7" => data <= "0000000000";
                when x"23F8" => data <= "0000000000";
                when x"23F9" => data <= "0000000000";
                when x"23FA" => data <= "0000000000";
                when x"23FB" => data <= "0000000000";
                when x"23FC" => data <= "0000000000";
                when x"23FD" => data <= "0000000000";
                when x"23FE" => data <= "0000000000";
                when x"23FF" => data <= "0000000000";
                when x"2400" => data <= "0000000000";
                when x"2401" => data <= "0000000000";
                when x"2402" => data <= "0000000000";
                when x"2403" => data <= "0000000000";
                when x"2404" => data <= "0000000000";
                when x"2405" => data <= "0000000000";
                when x"2406" => data <= "0000000000";
                when x"2407" => data <= "0000000000";
                when x"2408" => data <= "0000000000";
                when x"2409" => data <= "0000000000";
                when x"240A" => data <= "0000000000";
                when x"240B" => data <= "0000000000";
                when x"240C" => data <= "0000000000";
                when x"240D" => data <= "0000000000";
                when x"240E" => data <= "0000000000";
                when x"240F" => data <= "0000000000";
                when x"2410" => data <= "0000000000";
                when x"2411" => data <= "0000000000";
                when x"2412" => data <= "0000000000";
                when x"2413" => data <= "0000000000";
                when x"2414" => data <= "0000000000";
                when x"2415" => data <= "0000000000";
                when x"2416" => data <= "0000000000";
                when x"2417" => data <= "0000000000";
                when x"2418" => data <= "0000000000";
                when x"2419" => data <= "0000000000";
                when x"241A" => data <= "0000000000";
                when x"241B" => data <= "0000000000";
                when x"241C" => data <= "0000000000";
                when x"241D" => data <= "0000000000";
                when x"241E" => data <= "0000000000";
                when x"241F" => data <= "0000000000";
                when x"2420" => data <= "0000000000";
                when x"2421" => data <= "0000000000";
                when x"2422" => data <= "0000000000";
                when x"2423" => data <= "0000000000";
                when x"2424" => data <= "0000000000";
                when x"2425" => data <= "0000000000";
                when x"2426" => data <= "0000000000";
                when x"2427" => data <= "0000000000";
                when x"2428" => data <= "0000000000";
                when x"2429" => data <= "0000000000";
                when x"242A" => data <= "0000000000";
                when x"242B" => data <= "0000000000";
                when x"242C" => data <= "0000000000";
                when x"242D" => data <= "0000000000";
                when x"242E" => data <= "0000000000";
                when x"242F" => data <= "0000000000";
                when x"2430" => data <= "0000000000";
                when x"2431" => data <= "0000000000";
                when x"2432" => data <= "0000000000";
                when x"2433" => data <= "0000000000";
                when x"2434" => data <= "0000000000";
                when x"2435" => data <= "0000000000";
                when x"2436" => data <= "0000000000";
                when x"2437" => data <= "0000000000";
                when x"2438" => data <= "0000000000";
                when x"2439" => data <= "0000000000";
                when x"243A" => data <= "0000000000";
                when x"243B" => data <= "0000000000";
                when x"243C" => data <= "0000000000";
                when x"243D" => data <= "0000000000";
                when x"243E" => data <= "0000000000";
                when x"243F" => data <= "0000000000";
                when x"2440" => data <= "0000000000";
                when x"2441" => data <= "0000000000";
                when x"2442" => data <= "0000000000";
                when x"2443" => data <= "0000000000";
                when x"2444" => data <= "0000000000";
                when x"2445" => data <= "0000000000";
                when x"2446" => data <= "0000000000";
                when x"2447" => data <= "0000000000";
                when x"2448" => data <= "0000000000";
                when x"2449" => data <= "0000000000";
                when x"244A" => data <= "0000000000";
                when x"244B" => data <= "0000000000";
                when x"244C" => data <= "0000000000";
                when x"244D" => data <= "0000000000";
                when x"244E" => data <= "0000000000";
                when x"244F" => data <= "0000000000";
                when x"2450" => data <= "0000000000";
                when x"2451" => data <= "0000000000";
                when x"2452" => data <= "0000000000";
                when x"2453" => data <= "0000000000";
                when x"2454" => data <= "0000000000";
                when x"2455" => data <= "0000000000";
                when x"2456" => data <= "0000000000";
                when x"2457" => data <= "0000000000";
                when x"2458" => data <= "0000000000";
                when x"2459" => data <= "0000000000";
                when x"245A" => data <= "0000000000";
                when x"245B" => data <= "0000000000";
                when x"245C" => data <= "0000000000";
                when x"245D" => data <= "0000000000";
                when x"245E" => data <= "0000000000";
                when x"245F" => data <= "0000000000";
                when x"2460" => data <= "0000000000";
                when x"2461" => data <= "0000000000";
                when x"2462" => data <= "0000000000";
                when x"2463" => data <= "0000000000";
                when x"2464" => data <= "0000000000";
                when x"2465" => data <= "0000000000";
                when x"2466" => data <= "0000000000";
                when x"2467" => data <= "0000000000";
                when x"2468" => data <= "0000000000";
                when x"2469" => data <= "0000000000";
                when x"246A" => data <= "0000000000";
                when x"246B" => data <= "0000000000";
                when x"246C" => data <= "0000000000";
                when x"246D" => data <= "0000000000";
                when x"246E" => data <= "0000000000";
                when x"246F" => data <= "0000000000";
                when x"2470" => data <= "0000000000";
                when x"2471" => data <= "0000000000";
                when x"2472" => data <= "0000000000";
                when x"2473" => data <= "0000000000";
                when x"2474" => data <= "0000000000";
                when x"2475" => data <= "0000000000";
                when x"2476" => data <= "0110101000";
                when x"2477" => data <= "0000000000";
                when x"2478" => data <= "0000000000";
                when x"2479" => data <= "0000000000";
                when x"247A" => data <= "0000000000";
                when x"247B" => data <= "0000000000";
                when x"247C" => data <= "0000000000";
                when x"247D" => data <= "0000000000";
                when x"247E" => data <= "0000000000";
                when x"247F" => data <= "0000000000";
                when x"2480" => data <= "0000000000";
                when x"2481" => data <= "0000000000";
                when x"2482" => data <= "0000000000";
                when x"2483" => data <= "0000000000";
                when x"2484" => data <= "0000000000";
                when x"2485" => data <= "0000000000";
                when x"2486" => data <= "0000000000";
                when x"2487" => data <= "0000000000";
                when x"2488" => data <= "0000000000";
                when x"2489" => data <= "0000000000";
                when x"248A" => data <= "0000000000";
                when x"248B" => data <= "0000000000";
                when x"248C" => data <= "0000000000";
                when x"248D" => data <= "0000000000";
                when x"248E" => data <= "0000000000";
                when x"248F" => data <= "0000000000";
                when x"2490" => data <= "0000000000";
                when x"2491" => data <= "0000000000";
                when x"2492" => data <= "0000000000";
                when x"2493" => data <= "0000000000";
                when x"2494" => data <= "0000000000";
                when x"2495" => data <= "0000000000";
                when x"2496" => data <= "0000000000";
                when x"2497" => data <= "0000000000";
                when x"2498" => data <= "0000000000";
                when x"2499" => data <= "0000000000";
                when x"249A" => data <= "0000000000";
                when x"249B" => data <= "0000000000";
                when x"249C" => data <= "0000000000";
                when x"249D" => data <= "0000000000";
                when x"249E" => data <= "0000000000";
                when x"249F" => data <= "0000000000";
                when x"24A0" => data <= "0000000000";
                when x"24A1" => data <= "0000000000";
                when x"24A2" => data <= "0000000000";
                when x"24A3" => data <= "0000000000";
                when x"24A4" => data <= "0000000000";
                when x"24A5" => data <= "0000000000";
                when x"24A6" => data <= "0000000000";
                when x"24A7" => data <= "0000000000";
                when x"24A8" => data <= "0000000000";
                when x"24A9" => data <= "0000000000";
                when x"24AA" => data <= "0000000000";
                when x"24AB" => data <= "0000000000";
                when x"24AC" => data <= "0000000000";
                when x"24AD" => data <= "0000000000";
                when x"24AE" => data <= "0000000000";
                when x"24AF" => data <= "0000000000";
                when x"24B0" => data <= "0000000000";
                when x"24B1" => data <= "0000000000";
                when x"24B2" => data <= "0000000000";
                when x"24B3" => data <= "0000000000";
                when x"24B4" => data <= "0000000000";
                when x"24B5" => data <= "0000000000";
                when x"24B6" => data <= "0000000000";
                when x"24B7" => data <= "0000000000";
                when x"24B8" => data <= "0000000000";
                when x"24B9" => data <= "0000000000";
                when x"24BA" => data <= "0000000000";
                when x"24BB" => data <= "0000000000";
                when x"24BC" => data <= "0000000000";
                when x"24BD" => data <= "0000000000";
                when x"24BE" => data <= "0000000000";
                when x"24BF" => data <= "0000000000";
                when x"24C0" => data <= "0000000000";
                when x"24C1" => data <= "0000000000";
                when x"24C2" => data <= "0000000000";
                when x"24C3" => data <= "0000000000";
                when x"24C4" => data <= "0000000000";
                when x"24C5" => data <= "0000000000";
                when x"24C6" => data <= "0000000000";
                when x"24C7" => data <= "0000000000";
                when x"24C8" => data <= "0000000000";
                when x"24C9" => data <= "0000000000";
                when x"24CA" => data <= "0000000000";
                when x"24CB" => data <= "0000000000";
                when x"24CC" => data <= "0000000000";
                when x"24CD" => data <= "0000000000";
                when x"24CE" => data <= "0000000000";
                when x"24CF" => data <= "0000000000";
                when x"24D0" => data <= "0000000000";
                when x"24D1" => data <= "0000000000";
                when x"24D2" => data <= "0000000000";
                when x"24D3" => data <= "0000000000";
                when x"24D4" => data <= "0000000000";
                when x"24D5" => data <= "0000000000";
                when x"24D6" => data <= "0000000000";
                when x"24D7" => data <= "0000000000";
                when x"24D8" => data <= "0000000000";
                when x"24D9" => data <= "0000000000";
                when x"24DA" => data <= "0000000000";
                when x"24DB" => data <= "0000000000";
                when x"24DC" => data <= "0000000000";
                when x"24DD" => data <= "0000000000";
                when x"24DE" => data <= "0000000000";
                when x"24DF" => data <= "0000000000";
                when x"24E0" => data <= "0000000000";
                when x"24E1" => data <= "0000000000";
                when x"24E2" => data <= "0000000000";
                when x"24E3" => data <= "0000000000";
                when x"24E4" => data <= "0000000000";
                when x"24E5" => data <= "0000000000";
                when x"24E6" => data <= "0000000000";
                when x"24E7" => data <= "0000000000";
                when x"24E8" => data <= "0000000000";
                when x"24E9" => data <= "0000000000";
                when x"24EA" => data <= "0000000000";
                when x"24EB" => data <= "0000000000";
                when x"24EC" => data <= "0000000000";
                when x"24ED" => data <= "0000000000";
                when x"24EE" => data <= "0000000000";
                when x"24EF" => data <= "0000000000";
                when x"24F0" => data <= "0000000000";
                when x"24F1" => data <= "0000000000";
                when x"24F2" => data <= "0000000000";
                when x"24F3" => data <= "0000000000";
                when x"24F4" => data <= "0000000000";
                when x"24F5" => data <= "0000000000";
                when x"24F6" => data <= "0000000000";
                when x"24F7" => data <= "0000000000";
                when x"24F8" => data <= "0000000000";
                when x"24F9" => data <= "0000000000";
                when x"24FA" => data <= "0000000000";
                when x"24FB" => data <= "0000000000";
                when x"24FC" => data <= "0000000000";
                when x"24FD" => data <= "0000000000";
                when x"24FE" => data <= "0000000000";
                when x"24FF" => data <= "0000000000";
                when x"2500" => data <= "0000000000";
                when x"2501" => data <= "0000000000";
                when x"2502" => data <= "0000000000";
                when x"2503" => data <= "0000000000";
                when x"2504" => data <= "0000000000";
                when x"2505" => data <= "0000000000";
                when x"2506" => data <= "0000000000";
                when x"2507" => data <= "0000000000";
                when x"2508" => data <= "0000000000";
                when x"2509" => data <= "0000000000";
                when x"250A" => data <= "0000000000";
                when x"250B" => data <= "0000000000";
                when x"250C" => data <= "0000000000";
                when x"250D" => data <= "0000000000";
                when x"250E" => data <= "0000000000";
                when x"250F" => data <= "0000000000";
                when x"2510" => data <= "0000000000";
                when x"2511" => data <= "0000000000";
                when x"2512" => data <= "0000000000";
                when x"2513" => data <= "0000000000";
                when x"2514" => data <= "0000000000";
                when x"2515" => data <= "0000000000";
                when x"2516" => data <= "0000000000";
                when x"2517" => data <= "0000000000";
                when x"2518" => data <= "0000000000";
                when x"2519" => data <= "0000000000";
                when x"251A" => data <= "0000000000";
                when x"251B" => data <= "0000000000";
                when x"251C" => data <= "0000000000";
                when x"251D" => data <= "0000000000";
                when x"251E" => data <= "1001110011";
                when x"251F" => data <= "0000000000";
                when x"2520" => data <= "0000000000";
                when x"2521" => data <= "0000000000";
                when x"2522" => data <= "0000000000";
                when x"2523" => data <= "0000000000";
                when x"2524" => data <= "0000000000";
                when x"2525" => data <= "0000000000";
                when x"2526" => data <= "0000000000";
                when x"2527" => data <= "0000000000";
                when x"2528" => data <= "0000000000";
                when x"2529" => data <= "0000000000";
                when x"252A" => data <= "0000000000";
                when x"252B" => data <= "0000000000";
                when x"252C" => data <= "0000000000";
                when x"252D" => data <= "0000000000";
                when x"252E" => data <= "0000000000";
                when x"252F" => data <= "0000000000";
                when x"2530" => data <= "0000000000";
                when x"2531" => data <= "0000000000";
                when x"2532" => data <= "0000000000";
                when x"2533" => data <= "0000000000";
                when x"2534" => data <= "0000000000";
                when x"2535" => data <= "0000000000";
                when x"2536" => data <= "0000000000";
                when x"2537" => data <= "0000000000";
                when x"2538" => data <= "0000000000";
                when x"2539" => data <= "0000000000";
                when x"253A" => data <= "0000000000";
                when x"253B" => data <= "0000000000";
                when x"253C" => data <= "0000000000";
                when x"253D" => data <= "0000000000";
                when x"253E" => data <= "0000000000";
                when x"253F" => data <= "0000000000";
                when x"2540" => data <= "0000000000";
                when x"2541" => data <= "0000000000";
                when x"2542" => data <= "0000000000";
                when x"2543" => data <= "0000000000";
                when x"2544" => data <= "0000000000";
                when x"2545" => data <= "0000000000";
                when x"2546" => data <= "0000000000";
                when x"2547" => data <= "0000000000";
                when x"2548" => data <= "0000000000";
                when x"2549" => data <= "0000000000";
                when x"254A" => data <= "0000000000";
                when x"254B" => data <= "0000000000";
                when x"254C" => data <= "0000000000";
                when x"254D" => data <= "0000000000";
                when x"254E" => data <= "0000000000";
                when x"254F" => data <= "0000000000";
                when x"2550" => data <= "0000000000";
                when x"2551" => data <= "0000000000";
                when x"2552" => data <= "0000000000";
                when x"2553" => data <= "0000000000";
                when x"2554" => data <= "0000000000";
                when x"2555" => data <= "0000000000";
                when x"2556" => data <= "0000000000";
                when x"2557" => data <= "0000000000";
                when x"2558" => data <= "0000000000";
                when x"2559" => data <= "0000000000";
                when x"255A" => data <= "0000000000";
                when x"255B" => data <= "0000000000";
                when x"255C" => data <= "0000000000";
                when x"255D" => data <= "0000000000";
                when x"255E" => data <= "0000000000";
                when x"255F" => data <= "0000000000";
                when x"2560" => data <= "0000000000";
                when x"2561" => data <= "0000000000";
                when x"2562" => data <= "0000000000";
                when x"2563" => data <= "0000000000";
                when x"2564" => data <= "0000000000";
                when x"2565" => data <= "0000000000";
                when x"2566" => data <= "0000000000";
                when x"2567" => data <= "0000000000";
                when x"2568" => data <= "0000000000";
                when x"2569" => data <= "0000000000";
                when x"256A" => data <= "0000000000";
                when x"256B" => data <= "0000000000";
                when x"256C" => data <= "0000000000";
                when x"256D" => data <= "0000000000";
                when x"256E" => data <= "0000000000";
                when x"256F" => data <= "0000000000";
                when x"2570" => data <= "0000000000";
                when x"2571" => data <= "0000000000";
                when x"2572" => data <= "0000000000";
                when x"2573" => data <= "0000000000";
                when x"2574" => data <= "0000000000";
                when x"2575" => data <= "0111110111";
                when x"2576" => data <= "0000000000";
                when x"2577" => data <= "0000000000";
                when x"2578" => data <= "0000000000";
                when x"2579" => data <= "0000000000";
                when x"257A" => data <= "0000000000";
                when x"257B" => data <= "0000000000";
                when x"257C" => data <= "0000000000";
                when x"257D" => data <= "0000000000";
                when x"257E" => data <= "0000000000";
                when x"257F" => data <= "0000000000";
                when x"2580" => data <= "0000000000";
                when x"2581" => data <= "0000000000";
                when x"2582" => data <= "0000000000";
                when x"2583" => data <= "0000000000";
                when x"2584" => data <= "0000000000";
                when x"2585" => data <= "0000000000";
                when x"2586" => data <= "0000000000";
                when x"2587" => data <= "0000000000";
                when x"2588" => data <= "0000000000";
                when x"2589" => data <= "0000000000";
                when x"258A" => data <= "0000000000";
                when x"258B" => data <= "0000000000";
                when x"258C" => data <= "0000000000";
                when x"258D" => data <= "0000000000";
                when x"258E" => data <= "0000000000";
                when x"258F" => data <= "0000000000";
                when x"2590" => data <= "0000000000";
                when x"2591" => data <= "0000000000";
                when x"2592" => data <= "0000000000";
                when x"2593" => data <= "0000000000";
                when x"2594" => data <= "0000000000";
                when x"2595" => data <= "0000000000";
                when x"2596" => data <= "0000000000";
                when x"2597" => data <= "0000000000";
                when x"2598" => data <= "0000000000";
                when x"2599" => data <= "0000000000";
                when x"259A" => data <= "0000000000";
                when x"259B" => data <= "0000000000";
                when x"259C" => data <= "0000000000";
                when x"259D" => data <= "0000000000";
                when x"259E" => data <= "0000000000";
                when x"259F" => data <= "0000000000";
                when x"25A0" => data <= "0000000000";
                when x"25A1" => data <= "0000000000";
                when x"25A2" => data <= "0000000000";
                when x"25A3" => data <= "0000000000";
                when x"25A4" => data <= "0000000000";
                when x"25A5" => data <= "0000000000";
                when x"25A6" => data <= "0000000000";
                when x"25A7" => data <= "0000000000";
                when x"25A8" => data <= "0000000000";
                when x"25A9" => data <= "0000000000";
                when x"25AA" => data <= "0000000000";
                when x"25AB" => data <= "0000000000";
                when x"25AC" => data <= "0000000000";
                when x"25AD" => data <= "0000000000";
                when x"25AE" => data <= "0000000000";
                when x"25AF" => data <= "0000000000";
                when x"25B0" => data <= "0000000000";
                when x"25B1" => data <= "0000000000";
                when x"25B2" => data <= "0000000000";
                when x"25B3" => data <= "0000000000";
                when x"25B4" => data <= "0000000000";
                when x"25B5" => data <= "0000000000";
                when x"25B6" => data <= "0000000000";
                when x"25B7" => data <= "0000000000";
                when x"25B8" => data <= "0000000000";
                when x"25B9" => data <= "0000000000";
                when x"25BA" => data <= "0000000000";
                when x"25BB" => data <= "0000000000";
                when x"25BC" => data <= "0000000000";
                when x"25BD" => data <= "0000000000";
                when x"25BE" => data <= "0000000000";
                when x"25BF" => data <= "0000000000";
                when x"25C0" => data <= "0000000000";
                when x"25C1" => data <= "0000000000";
                when x"25C2" => data <= "0000000000";
                when x"25C3" => data <= "0000000000";
                when x"25C4" => data <= "0000000000";
                when x"25C5" => data <= "0000000000";
                when x"25C6" => data <= "0000000000";
                when x"25C7" => data <= "0000000000";
                when x"25C8" => data <= "0000000000";
                when x"25C9" => data <= "0000000000";
                when x"25CA" => data <= "0000000000";
                when x"25CB" => data <= "0000000000";
                when x"25CC" => data <= "0000000000";
                when x"25CD" => data <= "0000000000";
                when x"25CE" => data <= "0000000000";
                when x"25CF" => data <= "0000000000";
                when x"25D0" => data <= "0000000000";
                when x"25D1" => data <= "0000000000";
                when x"25D2" => data <= "0000000000";
                when x"25D3" => data <= "0000000000";
                when x"25D4" => data <= "0000000000";
                when x"25D5" => data <= "0000000000";
                when x"25D6" => data <= "0000000000";
                when x"25D7" => data <= "0000000000";
                when x"25D8" => data <= "0000000000";
                when x"25D9" => data <= "0000000000";
                when x"25DA" => data <= "0000000000";
                when x"25DB" => data <= "0000000000";
                when x"25DC" => data <= "0000000000";
                when x"25DD" => data <= "0000000000";
                when x"25DE" => data <= "0000000000";
                when x"25DF" => data <= "0000000000";
                when x"25E0" => data <= "0000000000";
                when x"25E1" => data <= "0000000000";
                when x"25E2" => data <= "0000000000";
                when x"25E3" => data <= "0000000000";
                when x"25E4" => data <= "0000000000";
                when x"25E5" => data <= "0000000000";
                when x"25E6" => data <= "0000000000";
                when x"25E7" => data <= "0000000000";
                when x"25E8" => data <= "0000000000";
                when x"25E9" => data <= "0000000000";
                when x"25EA" => data <= "0000000000";
                when x"25EB" => data <= "0000000000";
                when x"25EC" => data <= "0000000000";
                when x"25ED" => data <= "0000000000";
                when x"25EE" => data <= "0000000000";
                when x"25EF" => data <= "0000000000";
                when x"25F0" => data <= "0000000000";
                when x"25F1" => data <= "0000000000";
                when x"25F2" => data <= "0000000000";
                when x"25F3" => data <= "0000000000";
                when x"25F4" => data <= "0000000000";
                when x"25F5" => data <= "0000000000";
                when x"25F6" => data <= "0000000000";
                when x"25F7" => data <= "0000000000";
                when x"25F8" => data <= "0000000000";
                when x"25F9" => data <= "0000000000";
                when x"25FA" => data <= "0000000000";
                when x"25FB" => data <= "0000000000";
                when x"25FC" => data <= "0000000000";
                when x"25FD" => data <= "0000000000";
                when x"25FE" => data <= "0000000000";
                when x"25FF" => data <= "0000000000";
                when x"2600" => data <= "0000000000";
                when x"2601" => data <= "0000000000";
                when x"2602" => data <= "0000000000";
                when x"2603" => data <= "0000000000";
                when x"2604" => data <= "0111110111";
                when x"2605" => data <= "0000000000";
                when x"2606" => data <= "0000000000";
                when x"2607" => data <= "0000000000";
                when x"2608" => data <= "0000000000";
                when x"2609" => data <= "0000000000";
                when x"260A" => data <= "0000000000";
                when x"260B" => data <= "0000000000";
                when x"260C" => data <= "0000000000";
                when x"260D" => data <= "0000000000";
                when x"260E" => data <= "0000000000";
                when x"260F" => data <= "0000000000";
                when x"2610" => data <= "0000000000";
                when x"2611" => data <= "0000000000";
                when x"2612" => data <= "0000000000";
                when x"2613" => data <= "0000000000";
                when x"2614" => data <= "0000000000";
                when x"2615" => data <= "0000000000";
                when x"2616" => data <= "0000000000";
                when x"2617" => data <= "0000000000";
                when x"2618" => data <= "0000000000";
                when x"2619" => data <= "0000000000";
                when x"261A" => data <= "0000000000";
                when x"261B" => data <= "0000000000";
                when x"261C" => data <= "0000000000";
                when x"261D" => data <= "0000000000";
                when x"261E" => data <= "0000000000";
                when x"261F" => data <= "0000000000";
                when x"2620" => data <= "0000000000";
                when x"2621" => data <= "0000000000";
                when x"2622" => data <= "0000000000";
                when x"2623" => data <= "0000000000";
                when x"2624" => data <= "0000000000";
                when x"2625" => data <= "0000000000";
                when x"2626" => data <= "0000000000";
                when x"2627" => data <= "0000000000";
                when x"2628" => data <= "0000000000";
                when x"2629" => data <= "0000000000";
                when x"262A" => data <= "0000000000";
                when x"262B" => data <= "0000000000";
                when x"262C" => data <= "0000000000";
                when x"262D" => data <= "0000000000";
                when x"262E" => data <= "0000000000";
                when x"262F" => data <= "0000000000";
                when x"2630" => data <= "0000000000";
                when x"2631" => data <= "0000000000";
                when x"2632" => data <= "0000000000";
                when x"2633" => data <= "0000000000";
                when x"2634" => data <= "0000000000";
                when x"2635" => data <= "0000000000";
                when x"2636" => data <= "0000000000";
                when x"2637" => data <= "0000000000";
                when x"2638" => data <= "0000000000";
                when x"2639" => data <= "0000000000";
                when x"263A" => data <= "0000000000";
                when x"263B" => data <= "0000000000";
                when x"263C" => data <= "0000000000";
                when x"263D" => data <= "0000000000";
                when x"263E" => data <= "0000000000";
                when x"263F" => data <= "0000000000";
                when x"2640" => data <= "0000000000";
                when x"2641" => data <= "0000000000";
                when x"2642" => data <= "0000000000";
                when x"2643" => data <= "0000000000";
                when x"2644" => data <= "0000000000";
                when x"2645" => data <= "0000000000";
                when x"2646" => data <= "0000000000";
                when x"2647" => data <= "0000000000";
                when x"2648" => data <= "0000000000";
                when x"2649" => data <= "0000000000";
                when x"264A" => data <= "0000000000";
                when x"264B" => data <= "0000000000";
                when x"264C" => data <= "0000000000";
                when x"264D" => data <= "0000000000";
                when x"264E" => data <= "0000000000";
                when x"264F" => data <= "0000000000";
                when x"2650" => data <= "0000000000";
                when x"2651" => data <= "0000000000";
                when x"2652" => data <= "0000000000";
                when x"2653" => data <= "0000000000";
                when x"2654" => data <= "0000000000";
                when x"2655" => data <= "0000000000";
                when x"2656" => data <= "0000000000";
                when x"2657" => data <= "0000000000";
                when x"2658" => data <= "0000000000";
                when x"2659" => data <= "0000000000";
                when x"265A" => data <= "0000000000";
                when x"265B" => data <= "0000000000";
                when x"265C" => data <= "0000000000";
                when x"265D" => data <= "0000000000";
                when x"265E" => data <= "0000000000";
                when x"265F" => data <= "0000000000";
                when x"2660" => data <= "0000000000";
                when x"2661" => data <= "0000000000";
                when x"2662" => data <= "0000000000";
                when x"2663" => data <= "0000000000";
                when x"2664" => data <= "0000000000";
                when x"2665" => data <= "0000000000";
                when x"2666" => data <= "0000000000";
                when x"2667" => data <= "0000000000";
                when x"2668" => data <= "0000000000";
                when x"2669" => data <= "0000000000";
                when x"266A" => data <= "0000000000";
                when x"266B" => data <= "0000000000";
                when x"266C" => data <= "0000000000";
                when x"266D" => data <= "0000000000";
                when x"266E" => data <= "0000000000";
                when x"266F" => data <= "0000000000";
                when x"2670" => data <= "0000000000";
                when x"2671" => data <= "0111110111";
                when x"2672" => data <= "0000000000";
                when x"2673" => data <= "0000000000";
                when x"2674" => data <= "0000000000";
                when x"2675" => data <= "0000000000";
                when x"2676" => data <= "0000000000";
                when x"2677" => data <= "0000000000";
                when x"2678" => data <= "0000000000";
                when x"2679" => data <= "0000000000";
                when x"267A" => data <= "0000000000";
                when x"267B" => data <= "0000000000";
                when x"267C" => data <= "0000000000";
                when x"267D" => data <= "0000000000";
                when x"267E" => data <= "0000000000";
                when x"267F" => data <= "0000000000";
                when x"2680" => data <= "0000000000";
                when x"2681" => data <= "0000000000";
                when x"2682" => data <= "0000000000";
                when x"2683" => data <= "0000000000";
                when x"2684" => data <= "0000000000";
                when x"2685" => data <= "0000000000";
                when x"2686" => data <= "0000000000";
                when x"2687" => data <= "0000000000";
                when x"2688" => data <= "0000000000";
                when x"2689" => data <= "0000000000";
                when x"268A" => data <= "0000000000";
                when x"268B" => data <= "0000000000";
                when x"268C" => data <= "0000000000";
                when x"268D" => data <= "0000000000";
                when x"268E" => data <= "0000000000";
                when x"268F" => data <= "0000000000";
                when x"2690" => data <= "0000000000";
                when x"2691" => data <= "0000000000";
                when x"2692" => data <= "0000000000";
                when x"2693" => data <= "0000000000";
                when x"2694" => data <= "0000000000";
                when x"2695" => data <= "0000000000";
                when x"2696" => data <= "0000000000";
                when x"2697" => data <= "0000000000";
                when x"2698" => data <= "0000000000";
                when x"2699" => data <= "0000000000";
                when x"269A" => data <= "0000000000";
                when x"269B" => data <= "0000000000";
                when x"269C" => data <= "0000000000";
                when x"269D" => data <= "0000000000";
                when x"269E" => data <= "0000000000";
                when x"269F" => data <= "0000000000";
                when x"26A0" => data <= "0000000000";
                when x"26A1" => data <= "0000000000";
                when x"26A2" => data <= "0000000000";
                when x"26A3" => data <= "0000000000";
                when x"26A4" => data <= "0000000000";
                when x"26A5" => data <= "0000000000";
                when x"26A6" => data <= "0000000000";
                when x"26A7" => data <= "0000000000";
                when x"26A8" => data <= "0000000000";
                when x"26A9" => data <= "0000000000";
                when x"26AA" => data <= "0000000000";
                when x"26AB" => data <= "0000000000";
                when x"26AC" => data <= "0000000000";
                when x"26AD" => data <= "0000000000";
                when x"26AE" => data <= "0000000000";
                when x"26AF" => data <= "0000000000";
                when x"26B0" => data <= "0000000000";
                when x"26B1" => data <= "0000000000";
                when x"26B2" => data <= "0000000000";
                when x"26B3" => data <= "0000000000";
                when x"26B4" => data <= "0000000000";
                when x"26B5" => data <= "0000000000";
                when x"26B6" => data <= "0000000000";
                when x"26B7" => data <= "0000000000";
                when x"26B8" => data <= "0000000000";
                when x"26B9" => data <= "0000000000";
                when x"26BA" => data <= "0000000000";
                when x"26BB" => data <= "0000000000";
                when x"26BC" => data <= "0000000000";
                when x"26BD" => data <= "0000000000";
                when x"26BE" => data <= "0000000000";
                when x"26BF" => data <= "0000000000";
                when x"26C0" => data <= "0000000000";
                when x"26C1" => data <= "0000000000";
                when x"26C2" => data <= "0000000000";
                when x"26C3" => data <= "0000000000";
                when x"26C4" => data <= "0000000000";
                when x"26C5" => data <= "0000000000";
                when x"26C6" => data <= "0000000000";
                when x"26C7" => data <= "0000000000";
                when x"26C8" => data <= "0000000000";
                when x"26C9" => data <= "0000000000";
                when x"26CA" => data <= "0000000000";
                when x"26CB" => data <= "0000000000";
                when x"26CC" => data <= "0000000000";
                when x"26CD" => data <= "0000000000";
                when x"26CE" => data <= "0000000000";
                when x"26CF" => data <= "0000000000";
                when x"26D0" => data <= "0000000000";
                when x"26D1" => data <= "0000000000";
                when x"26D2" => data <= "0000000000";
                when x"26D3" => data <= "0000000000";
                when x"26D4" => data <= "0000000000";
                when x"26D5" => data <= "0000000000";
                when x"26D6" => data <= "0000000000";
                when x"26D7" => data <= "0000000000";
                when x"26D8" => data <= "0000000000";
                when x"26D9" => data <= "0000000000";
                when x"26DA" => data <= "0000000000";
                when x"26DB" => data <= "0000000000";
                when x"26DC" => data <= "0000000000";
                when x"26DD" => data <= "0000000000";
                when x"26DE" => data <= "0000000000";
                when x"26DF" => data <= "0000000000";
                when x"26E0" => data <= "0000000000";
                when x"26E1" => data <= "0000000000";
                when x"26E2" => data <= "0000000000";
                when x"26E3" => data <= "0000000000";
                when x"26E4" => data <= "0000000000";
                when x"26E5" => data <= "0000000000";
                when x"26E6" => data <= "0000000000";
                when x"26E7" => data <= "0000000000";
                when x"26E8" => data <= "0000000000";
                when x"26E9" => data <= "0000000000";
                when x"26EA" => data <= "0000000000";
                when x"26EB" => data <= "0000000000";
                when x"26EC" => data <= "0000000000";
                when x"26ED" => data <= "0000000000";
                when x"26EE" => data <= "0000000000";
                when x"26EF" => data <= "0000000000";
                when x"26F0" => data <= "0000000000";
                when x"26F1" => data <= "0000000000";
                when x"26F2" => data <= "0000000000";
                when x"26F3" => data <= "0000000000";
                when x"26F4" => data <= "0000000000";
                when x"26F5" => data <= "0000000000";
                when x"26F6" => data <= "0000000000";
                when x"26F7" => data <= "0000000000";
                when x"26F8" => data <= "0000000000";
                when x"26F9" => data <= "0000000000";
                when x"26FA" => data <= "0000000000";
                when x"26FB" => data <= "0000000000";
                when x"26FC" => data <= "0000000000";
                when x"26FD" => data <= "0000000000";
                when x"26FE" => data <= "0000000000";
                when x"26FF" => data <= "0000000000";
                when x"2700" => data <= "0000000000";
                when x"2701" => data <= "0000000000";
                when x"2702" => data <= "0000000000";
                when x"2703" => data <= "0000000000";
                when x"2704" => data <= "0000000000";
                when x"2705" => data <= "0000000000";
                when x"2706" => data <= "0000000000";
                when x"2707" => data <= "0000000000";
                when x"2708" => data <= "0000000000";
                when x"2709" => data <= "0000000000";
                when x"270A" => data <= "0000000000";
                when x"270B" => data <= "0000000000";
                when x"270C" => data <= "0000000000";
                when x"270D" => data <= "0000000000";
                when x"270E" => data <= "0000000000";
                when x"270F" => data <= "0000000000";
                when x"2710" => data <= "0000000000";
                when x"2711" => data <= "0000000000";
                when x"2712" => data <= "0000000000";
                when x"2713" => data <= "0000000000";
                when x"2714" => data <= "0000000000";
                when x"2715" => data <= "0000000000";
                when x"2716" => data <= "0000000000";
                when x"2717" => data <= "0000000000";
                when x"2718" => data <= "0000000000";
                when x"2719" => data <= "0000000000";
                when x"271A" => data <= "0000000000";
                when x"271B" => data <= "0000000000";
                when x"271C" => data <= "0000000000";
                when x"271D" => data <= "0000000000";
                when x"271E" => data <= "0000000000";
                when x"271F" => data <= "0000000000";
                when x"2720" => data <= "0000000000";
                when x"2721" => data <= "0000000000";
                when x"2722" => data <= "0000000000";
                when x"2723" => data <= "0000000000";
                when x"2724" => data <= "0000000000";
                when x"2725" => data <= "0000000000";
                when x"2726" => data <= "0000000000";
                when x"2727" => data <= "0000000000";
                when x"2728" => data <= "0000000000";
                when x"2729" => data <= "0000000000";
                when x"272A" => data <= "0000000000";
                when x"272B" => data <= "0000000000";
                when x"272C" => data <= "0000000000";
                when x"272D" => data <= "0000000000";
                when x"272E" => data <= "0000000000";
                when x"272F" => data <= "0000000000";
                when x"2730" => data <= "0000000000";
                when x"2731" => data <= "0000000000";
                when x"2732" => data <= "0000000000";
                when x"2733" => data <= "0000000000";
                when x"2734" => data <= "0000000000";
                when x"2735" => data <= "0000000000";
                when x"2736" => data <= "0000000000";
                when x"2737" => data <= "0000000000";
                when x"2738" => data <= "0000000000";
                when x"2739" => data <= "0000000000";
                when x"273A" => data <= "0000000000";
                when x"273B" => data <= "0000000000";
                when x"273C" => data <= "0000000000";
                when x"273D" => data <= "0000000000";
                when x"273E" => data <= "0000000000";
                when x"273F" => data <= "0000000000";
                when x"2740" => data <= "0000000000";
                when x"2741" => data <= "0000000000";
                when x"2742" => data <= "0000000000";
                when x"2743" => data <= "0000000000";
                when x"2744" => data <= "0000000000";
                when x"2745" => data <= "0000000000";
                when x"2746" => data <= "0000000000";
                when x"2747" => data <= "0000000000";
                when x"2748" => data <= "0000000000";
                when x"2749" => data <= "0000000000";
                when x"274A" => data <= "0000000000";
                when x"274B" => data <= "0000000000";
                when x"274C" => data <= "0000000000";
                when x"274D" => data <= "0000000000";
                when x"274E" => data <= "0000000000";
                when x"274F" => data <= "0000000000";
                when x"2750" => data <= "0000000000";
                when x"2751" => data <= "0000000000";
                when x"2752" => data <= "0000000000";
                when x"2753" => data <= "0000000000";
                when x"2754" => data <= "0000000000";
                when x"2755" => data <= "0000000000";
                when x"2756" => data <= "0000000000";
                when x"2757" => data <= "0000000000";
                when x"2758" => data <= "0000000000";
                when x"2759" => data <= "0000000000";
                when x"275A" => data <= "0000000000";
                when x"275B" => data <= "0000000000";
                when x"275C" => data <= "0000000000";
                when x"275D" => data <= "0000000000";
                when x"275E" => data <= "0000000000";
                when x"275F" => data <= "0000000000";
                when x"2760" => data <= "0000000000";
                when x"2761" => data <= "0000000000";
                when x"2762" => data <= "0000000000";
                when x"2763" => data <= "0000000000";
                when x"2764" => data <= "0000000000";
                when x"2765" => data <= "0000000000";
                when x"2766" => data <= "0000000000";
                when x"2767" => data <= "0000000000";
                when x"2768" => data <= "0000000000";
                when x"2769" => data <= "0000000000";
                when x"276A" => data <= "0000000000";
                when x"276B" => data <= "0000000000";
                when x"276C" => data <= "0000000000";
                when x"276D" => data <= "0000000000";
                when x"276E" => data <= "0000000000";
                when x"276F" => data <= "0000000000";
                when x"2770" => data <= "0000000000";
                when x"2771" => data <= "0000000000";
                when x"2772" => data <= "0000000000";
                when x"2773" => data <= "0000000000";
                when x"2774" => data <= "0000000000";
                when x"2775" => data <= "0000000000";
                when x"2776" => data <= "0000000000";
                when x"2777" => data <= "0000000000";
                when x"2778" => data <= "0000000000";
                when x"2779" => data <= "0000000000";
                when x"277A" => data <= "0000000000";
                when x"277B" => data <= "0000000000";
                when x"277C" => data <= "0000000000";
                when x"277D" => data <= "0000000000";
                when x"277E" => data <= "0000000000";
                when x"277F" => data <= "0000000000";
                when x"2780" => data <= "0000000000";
                when x"2781" => data <= "0000000000";
                when x"2782" => data <= "0000000000";
                when x"2783" => data <= "0000000000";
                when x"2784" => data <= "0000000000";
                when x"2785" => data <= "0000000000";
                when x"2786" => data <= "0000000000";
                when x"2787" => data <= "0000000000";
                when x"2788" => data <= "0000000000";
                when x"2789" => data <= "0000000000";
                when x"278A" => data <= "0000000000";
                when x"278B" => data <= "0000000000";
                when x"278C" => data <= "0000000000";
                when x"278D" => data <= "0000000000";
                when x"278E" => data <= "0000000000";
                when x"278F" => data <= "0000000000";
                when x"2790" => data <= "0000000000";
                when x"2791" => data <= "0000000000";
                when x"2792" => data <= "0000000000";
                when x"2793" => data <= "0000000000";
                when x"2794" => data <= "0000000000";
                when x"2795" => data <= "0000000000";
                when x"2796" => data <= "0000000000";
                when x"2797" => data <= "0000000000";
                when x"2798" => data <= "0000000000";
                when x"2799" => data <= "0000000000";
                when x"279A" => data <= "0000000000";
                when x"279B" => data <= "0000000000";
                when x"279C" => data <= "0000000000";
                when x"279D" => data <= "0000000000";
                when x"279E" => data <= "0000000000";
                when x"279F" => data <= "0000000000";
                when x"27A0" => data <= "0000000000";
                when x"27A1" => data <= "0000000000";
                when x"27A2" => data <= "0000000000";
                when x"27A3" => data <= "0000000000";
                when x"27A4" => data <= "0000000000";
                when x"27A5" => data <= "0000000000";
                when x"27A6" => data <= "0000000000";
                when x"27A7" => data <= "0000000000";
                when x"27A8" => data <= "0000000000";
                when x"27A9" => data <= "0000000000";
                when x"27AA" => data <= "0000000000";
                when x"27AB" => data <= "0000000000";
                when x"27AC" => data <= "0000000000";
                when x"27AD" => data <= "0000000000";
                when x"27AE" => data <= "0000000000";
                when x"27AF" => data <= "0000000000";
                when x"27B0" => data <= "0000000000";
                when x"27B1" => data <= "0000000000";
                when x"27B2" => data <= "0000000000";
                when x"27B3" => data <= "0000000000";
                when x"27B4" => data <= "0000000000";
                when x"27B5" => data <= "0000000000";
                when x"27B6" => data <= "0000000000";
                when x"27B7" => data <= "0000000000";
                when x"27B8" => data <= "0000000000";
                when x"27B9" => data <= "0000000000";
                when x"27BA" => data <= "0000000000";
                when x"27BB" => data <= "0000000000";
                when x"27BC" => data <= "0000000000";
                when x"27BD" => data <= "0000000000";
                when x"27BE" => data <= "0000000000";
                when x"27BF" => data <= "0000000000";
                when x"27C0" => data <= "0000000000";
                when x"27C1" => data <= "0000000000";
                when x"27C2" => data <= "0000000000";
                when x"27C3" => data <= "0000000000";
                when x"27C4" => data <= "0000000000";
                when x"27C5" => data <= "0000000000";
                when x"27C6" => data <= "0000000000";
                when x"27C7" => data <= "0000000000";
                when x"27C8" => data <= "0000000000";
                when x"27C9" => data <= "0000000000";
                when x"27CA" => data <= "0000000000";
                when x"27CB" => data <= "0000000000";
                when x"27CC" => data <= "0000000000";
                when x"27CD" => data <= "0000000000";
                when x"27CE" => data <= "0000000000";
                when x"27CF" => data <= "0000000000";
                when x"27D0" => data <= "0000000000";
                when x"27D1" => data <= "0000000000";
                when x"27D2" => data <= "0000000000";
                when x"27D3" => data <= "0000000000";
                when x"27D4" => data <= "0000000000";
                when x"27D5" => data <= "0000000000";
                when x"27D6" => data <= "0000000000";
                when x"27D7" => data <= "0000000000";
                when x"27D8" => data <= "0000000000";
                when x"27D9" => data <= "0000000000";
                when x"27DA" => data <= "0000000000";
                when x"27DB" => data <= "0000000000";
                when x"27DC" => data <= "0000000000";
                when x"27DD" => data <= "0000000000";
                when x"27DE" => data <= "0000000000";
                when x"27DF" => data <= "0000000000";
                when x"27E0" => data <= "0000000000";
                when x"27E1" => data <= "0000000000";
                when x"27E2" => data <= "0000000000";
                when x"27E3" => data <= "0000000000";
                when x"27E4" => data <= "0000000000";
                when x"27E5" => data <= "0000000000";
                when x"27E6" => data <= "0000000000";
                when x"27E7" => data <= "0000000000";
                when x"27E8" => data <= "0000000000";
                when x"27E9" => data <= "0000000000";
                when x"27EA" => data <= "0000000000";
                when x"27EB" => data <= "0000000000";
                when x"27EC" => data <= "0000000000";
                when x"27ED" => data <= "0000000000";
                when x"27EE" => data <= "0000000000";
                when x"27EF" => data <= "0000000000";
                when x"27F0" => data <= "0000000000";
                when x"27F1" => data <= "0000000000";
                when x"27F2" => data <= "0000000000";
                when x"27F3" => data <= "0000000000";
                when x"27F4" => data <= "0000000000";
                when x"27F5" => data <= "0000000000";
                when x"27F6" => data <= "0000000000";
                when x"27F7" => data <= "0000000000";
                when x"27F8" => data <= "0000000000";
                when x"27F9" => data <= "0000000000";
                when x"27FA" => data <= "0000000000";
                when x"27FB" => data <= "0000000000";
                when x"27FC" => data <= "0000000000";
                when x"27FD" => data <= "0000000000";
                when x"27FE" => data <= "0000000000";
                when x"27FF" => data <= "0000000000";
                when others => data <= (others => '0');
            end case;
        end if;
    end process;
end Behavioral;

------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ECC_CHV_img_10000 is
    Port (
        clk     : in  STD_LOGIC;
        address : in  STD_LOGIC_VECTOR(13 downto 0);
        data    : out STD_LOGIC_VECTOR(5 downto 0)
    );
end ECC_CHV_img_10000;

architecture Behavioral of ECC_CHV_img_10000 is
begin
    process(clk)
    begin
        if rising_edge(clk) then
            case address is
                when x"00" => data <= "00000";
                when x"01" => data <= "00000";
                when x"02" => data <= "00000";
                when x"03" => data <= "00000";
                when x"04" => data <= "00000";
                when x"05" => data <= "00000";
                when x"06" => data <= "00000";
                when x"07" => data <= "00000";
                when x"08" => data <= "00000";
                when x"09" => data <= "00000";
                when x"0A" => data <= "00000";
                when x"0B" => data <= "00000";
                when x"0C" => data <= "00000";
                when x"0D" => data <= "00000";
                when x"0E" => data <= "00000";
                when x"0F" => data <= "00000";
                when x"10" => data <= "00000";
                when x"11" => data <= "00000";
                when x"12" => data <= "00000";
                when x"13" => data <= "00000";
                when x"14" => data <= "00000";
                when x"15" => data <= "00000";
                when x"16" => data <= "00000";
                when x"17" => data <= "00000";
                when x"18" => data <= "00000";
                when x"19" => data <= "00000";
                when x"1A" => data <= "00000";
                when x"1B" => data <= "00000";
                when x"1C" => data <= "00000";
                when x"1D" => data <= "00000";
                when x"1E" => data <= "00000";
                when x"1F" => data <= "00000";
                when x"20" => data <= "00000";
                when x"21" => data <= "00000";
                when x"22" => data <= "00000";
                when x"23" => data <= "00000";
                when x"24" => data <= "00000";
                when x"25" => data <= "00000";
                when x"26" => data <= "00000";
                when x"27" => data <= "00000";
                when x"28" => data <= "00000";
                when x"29" => data <= "00000";
                when x"2A" => data <= "00000";
                when x"2B" => data <= "00000";
                when x"2C" => data <= "00000";
                when x"2D" => data <= "00000";
                when x"2E" => data <= "00000";
                when x"2F" => data <= "00000";
                when x"30" => data <= "00000";
                when x"31" => data <= "00000";
                when x"32" => data <= "00000";
                when x"33" => data <= "00000";
                when x"34" => data <= "00000";
                when x"35" => data <= "00000";
                when x"36" => data <= "00000";
                when x"37" => data <= "00000";
                when x"38" => data <= "00000";
                when x"39" => data <= "00000";
                when x"3A" => data <= "00000";
                when x"3B" => data <= "00000";
                when x"3C" => data <= "00000";
                when x"3D" => data <= "00000";
                when x"3E" => data <= "00000";
                when x"3F" => data <= "00000";
                when x"40" => data <= "00000";
                when x"41" => data <= "00000";
                when x"42" => data <= "00000";
                when x"43" => data <= "00000";
                when x"44" => data <= "00000";
                when x"45" => data <= "00000";
                when x"46" => data <= "00000";
                when x"47" => data <= "00000";
                when x"48" => data <= "00000";
                when x"49" => data <= "00000";
                when x"4A" => data <= "00000";
                when x"4B" => data <= "00000";
                when x"4C" => data <= "00000";
                when x"4D" => data <= "00000";
                when x"4E" => data <= "00000";
                when x"4F" => data <= "00000";
                when x"50" => data <= "00000";
                when x"51" => data <= "00000";
                when x"52" => data <= "00000";
                when x"53" => data <= "00000";
                when x"54" => data <= "00000";
                when x"55" => data <= "00000";
                when x"56" => data <= "00000";
                when x"57" => data <= "00000";
                when x"58" => data <= "00000";
                when x"59" => data <= "00000";
                when x"5A" => data <= "00000";
                when x"5B" => data <= "00000";
                when x"5C" => data <= "00000";
                when x"5D" => data <= "00000";
                when x"5E" => data <= "00000";
                when x"5F" => data <= "00000";
                when x"60" => data <= "00000";
                when x"61" => data <= "00000";
                when x"62" => data <= "00000";
                when x"63" => data <= "00000";
                when x"64" => data <= "00000";
                when x"65" => data <= "00000";
                when x"66" => data <= "00000";
                when x"67" => data <= "00000";
                when x"68" => data <= "00000";
                when x"69" => data <= "00000";
                when x"6A" => data <= "00000";
                when x"6B" => data <= "00000";
                when x"6C" => data <= "00000";
                when x"6D" => data <= "00000";
                when x"6E" => data <= "00000";
                when x"6F" => data <= "00000";
                when x"70" => data <= "00000";
                when x"71" => data <= "00000";
                when x"72" => data <= "00000";
                when x"73" => data <= "00000";
                when x"74" => data <= "00000";
                when x"75" => data <= "00000";
                when x"76" => data <= "00000";
                when x"77" => data <= "00000";
                when x"78" => data <= "00000";
                when x"79" => data <= "00000";
                when x"7A" => data <= "00000";
                when x"7B" => data <= "00000";
                when x"7C" => data <= "00000";
                when x"7D" => data <= "00000";
                when x"7E" => data <= "00000";
                when x"7F" => data <= "00000";
                when x"80" => data <= "00000";
                when x"81" => data <= "00000";
                when x"82" => data <= "00000";
                when x"83" => data <= "00000";
                when x"84" => data <= "00000";
                when x"85" => data <= "00000";
                when x"86" => data <= "00000";
                when x"87" => data <= "00000";
                when x"88" => data <= "00000";
                when x"89" => data <= "00000";
                when x"8A" => data <= "00000";
                when x"8B" => data <= "00000";
                when x"8C" => data <= "00000";
                when x"8D" => data <= "00000";
                when x"8E" => data <= "00000";
                when x"8F" => data <= "00000";
                when x"90" => data <= "00000";
                when x"91" => data <= "00000";
                when x"92" => data <= "00000";
                when x"93" => data <= "00000";
                when x"94" => data <= "00000";
                when x"95" => data <= "00000";
                when x"96" => data <= "00000";
                when x"97" => data <= "00000";
                when x"98" => data <= "00000";
                when x"99" => data <= "00000";
                when x"9A" => data <= "00000";
                when x"9B" => data <= "00000";
                when x"9C" => data <= "00000";
                when x"9D" => data <= "00000";
                when x"9E" => data <= "00000";
                when x"9F" => data <= "00000";
                when x"A0" => data <= "00000";
                when x"A1" => data <= "00000";
                when x"A2" => data <= "00000";
                when x"A3" => data <= "00000";
                when x"A4" => data <= "00000";
                when x"A5" => data <= "00000";
                when x"A6" => data <= "00000";
                when x"A7" => data <= "00000";
                when x"A8" => data <= "00000";
                when x"A9" => data <= "00000";
                when x"AA" => data <= "00000";
                when x"AB" => data <= "00000";
                when x"AC" => data <= "00000";
                when x"AD" => data <= "00000";
                when x"AE" => data <= "00000";
                when x"AF" => data <= "00000";
                when x"B0" => data <= "00000";
                when x"B1" => data <= "00000";
                when x"B2" => data <= "00000";
                when x"B3" => data <= "00000";
                when x"B4" => data <= "00000";
                when x"B5" => data <= "00000";
                when x"B6" => data <= "00000";
                when x"B7" => data <= "00000";
                when x"B8" => data <= "00000";
                when x"B9" => data <= "00000";
                when x"BA" => data <= "00000";
                when x"BB" => data <= "00000";
                when x"BC" => data <= "00000";
                when x"BD" => data <= "00000";
                when x"BE" => data <= "00000";
                when x"BF" => data <= "00000";
                when x"C0" => data <= "00000";
                when x"C1" => data <= "00000";
                when x"C2" => data <= "00000";
                when x"C3" => data <= "00000";
                when x"C4" => data <= "00000";
                when x"C5" => data <= "00000";
                when x"C6" => data <= "00000";
                when x"C7" => data <= "00000";
                when x"C8" => data <= "00000";
                when x"C9" => data <= "00000";
                when x"CA" => data <= "00000";
                when x"CB" => data <= "00000";
                when x"CC" => data <= "00000";
                when x"CD" => data <= "00000";
                when x"CE" => data <= "00000";
                when x"CF" => data <= "00000";
                when x"D0" => data <= "00000";
                when x"D1" => data <= "00000";
                when x"D2" => data <= "00000";
                when x"D3" => data <= "00000";
                when x"D4" => data <= "00000";
                when x"D5" => data <= "00000";
                when x"D6" => data <= "00000";
                when x"D7" => data <= "00000";
                when x"D8" => data <= "00000";
                when x"D9" => data <= "00000";
                when x"DA" => data <= "00000";
                when x"DB" => data <= "00000";
                when x"DC" => data <= "00000";
                when x"DD" => data <= "00000";
                when x"DE" => data <= "00000";
                when x"DF" => data <= "00000";
                when x"E0" => data <= "00000";
                when x"E1" => data <= "00000";
                when x"E2" => data <= "00000";
                when x"E3" => data <= "00000";
                when x"E4" => data <= "00000";
                when x"E5" => data <= "00000";
                when x"E6" => data <= "00000";
                when x"E7" => data <= "00000";
                when x"E8" => data <= "00000";
                when x"E9" => data <= "00000";
                when x"EA" => data <= "00000";
                when x"EB" => data <= "00000";
                when x"EC" => data <= "00000";
                when x"ED" => data <= "00000";
                when x"EE" => data <= "00000";
                when x"EF" => data <= "00000";
                when x"F0" => data <= "00011";
                when x"F1" => data <= "00110";
                when x"F2" => data <= "00110";
                when x"F3" => data <= "11011";
                when x"F4" => data <= "00110";
                when x"F5" => data <= "00110";
                when x"F6" => data <= "00000";
                when x"F7" => data <= "00110";
                when x"F8" => data <= "00000";
                when x"F9" => data <= "01101";
                when x"FA" => data <= "00000";
                when x"FB" => data <= "00000";
                when x"FC" => data <= "00000";
                when x"FD" => data <= "00110";
                when x"FE" => data <= "00110";
                when x"FF" => data <= "00110";
                when x"100" => data <= "00110";
                when x"101" => data <= "10010";
                when x"102" => data <= "00000";
                when x"103" => data <= "00000";
                when x"104" => data <= "01011";
                when x"105" => data <= "01011";
                when x"106" => data <= "00000";
                when x"107" => data <= "00110";
                when x"108" => data <= "00110";
                when x"109" => data <= "00000";
                when x"10A" => data <= "00000";
                when x"10B" => data <= "00110";
                when x"10C" => data <= "01011";
                when x"10D" => data <= "00110";
                when x"10E" => data <= "00110";
                when x"10F" => data <= "10101";
                when x"110" => data <= "00110";
                when x"111" => data <= "00110";
                when x"112" => data <= "00110";
                when x"113" => data <= "00110";
                when x"114" => data <= "00110";
                when x"115" => data <= "00000";
                when x"116" => data <= "00110";
                when x"117" => data <= "00000";
                when x"118" => data <= "11111";
                when x"119" => data <= "00000";
                when x"11A" => data <= "11010";
                when x"11B" => data <= "01011";
                when x"11C" => data <= "00000";
                when x"11D" => data <= "00110";
                when x"11E" => data <= "10111";
                when x"11F" => data <= "00110";
                when x"120" => data <= "00010";
                when x"121" => data <= "00110";
                when x"122" => data <= "10011";
                when x"123" => data <= "01100";
                when x"124" => data <= "01011";
                when x"125" => data <= "00110";
                when x"126" => data <= "00000";
                when x"127" => data <= "10001";
                when x"128" => data <= "00110";
                when x"129" => data <= "00110";
                when x"12A" => data <= "00110";
                when x"12B" => data <= "00000";
                when x"12C" => data <= "00110";
                when x"12D" => data <= "00110";
                when x"12E" => data <= "00110";
                when x"12F" => data <= "00110";
                when x"130" => data <= "01101";
                when x"131" => data <= "00000";
                when x"132" => data <= "00110";
                when x"133" => data <= "00000";
                when x"134" => data <= "00110";
                when x"135" => data <= "00110";
                when x"136" => data <= "00110";
                when x"137" => data <= "11001";
                when x"138" => data <= "00110";
                when x"139" => data <= "00000";
                when x"13A" => data <= "11111";
                when x"13B" => data <= "00110";
                when x"13C" => data <= "00110";
                when x"13D" => data <= "00110";
                when x"13E" => data <= "00000";
                when x"13F" => data <= "01101";
                when x"140" => data <= "10011";
                when x"141" => data <= "00110";
                when x"142" => data <= "11001";
                when x"143" => data <= "00000";
                when x"144" => data <= "00000";
                when x"145" => data <= "00000";
                when x"146" => data <= "10001";
                when x"147" => data <= "00000";
                when x"148" => data <= "00001";
                when x"149" => data <= "00000";
                when x"14A" => data <= "00000";
                when x"14B" => data <= "10101";
                when x"14C" => data <= "00000";
                when x"14D" => data <= "00110";
                when x"14E" => data <= "11000";
                when x"14F" => data <= "00110";
                when x"150" => data <= "00000";
                when x"151" => data <= "00110";
                when x"152" => data <= "00110";
                when x"153" => data <= "00110";
                when x"154" => data <= "00110";
                when x"155" => data <= "00110";
                when x"156" => data <= "00110";
                when x"157" => data <= "00000";
                when x"158" => data <= "00000";
                when x"159" => data <= "00000";
                when x"15A" => data <= "00110";
                when x"15B" => data <= "01101";
                when x"15C" => data <= "00110";
                when x"15D" => data <= "11001";
                when x"15E" => data <= "00101";
                when x"15F" => data <= "00110";
                when x"160" => data <= "00101";
                when x"161" => data <= "00000";
                when x"162" => data <= "00000";
                when x"163" => data <= "00000";
                when x"164" => data <= "11100";
                when x"165" => data <= "00110";
                when x"166" => data <= "00110";
                when x"167" => data <= "00000";
                when x"168" => data <= "00000";
                when x"169" => data <= "10000";
                when x"16A" => data <= "10010";
                when x"16B" => data <= "00110";
                when x"16C" => data <= "00111";
                when x"16D" => data <= "00110";
                when x"16E" => data <= "00110";
                when x"16F" => data <= "00000";
                when x"170" => data <= "00001";
                when x"171" => data <= "00000";
                when x"172" => data <= "00000";
                when x"173" => data <= "00000";
                when x"174" => data <= "10010";
                when x"175" => data <= "00110";
                when x"176" => data <= "00110";
                when x"177" => data <= "00110";
                when x"178" => data <= "00110";
                when x"179" => data <= "00110";
                when x"17A" => data <= "11111";
                when x"17B" => data <= "01110";
                when x"17C" => data <= "00110";
                when x"17D" => data <= "00000";
                when x"17E" => data <= "00110";
                when x"17F" => data <= "00110";
                when x"180" => data <= "00000";
                when x"181" => data <= "00110";
                when x"182" => data <= "00110";
                when x"183" => data <= "01101";
                when x"184" => data <= "00000";
                when x"185" => data <= "00000";
                when x"186" => data <= "00110";
                when x"187" => data <= "10101";
                when x"188" => data <= "00110";
                when x"189" => data <= "00000";
                when x"18A" => data <= "00000";
                when x"18B" => data <= "00110";
                when x"18C" => data <= "00000";
                when x"18D" => data <= "00110";
                when x"18E" => data <= "00110";
                when x"18F" => data <= "00000";
                when x"190" => data <= "00000";
                when x"191" => data <= "00110";
                when x"192" => data <= "00110";
                when x"193" => data <= "00110";
                when x"194" => data <= "00110";
                when x"195" => data <= "00000";
                when x"196" => data <= "00000";
                when x"197" => data <= "00110";
                when x"198" => data <= "00000";
                when x"199" => data <= "00000";
                when x"19A" => data <= "00110";
                when x"19B" => data <= "00000";
                when x"19C" => data <= "00000";
                when x"19D" => data <= "00000";
                when x"19E" => data <= "01111";
                when x"19F" => data <= "00110";
                when x"1A0" => data <= "00110";
                when x"1A1" => data <= "01011";
                when x"1A2" => data <= "00110";
                when x"1A3" => data <= "00000";
                when x"1A4" => data <= "00000";
                when x"1A5" => data <= "00110";
                when x"1A6" => data <= "00110";
                when x"1A7" => data <= "00000";
                when x"1A8" => data <= "01010";
                when x"1A9" => data <= "00110";
                when x"1AA" => data <= "00000";
                when x"1AB" => data <= "00110";
                when x"1AC" => data <= "11000";
                when x"1AD" => data <= "00000";
                when x"1AE" => data <= "00110";
                when x"1AF" => data <= "00110";
                when x"1B0" => data <= "00000";
                when x"1B1" => data <= "00000";
                when x"1B2" => data <= "00000";
                when x"1B3" => data <= "00000";
                when x"1B4" => data <= "00110";
                when x"1B5" => data <= "11100";
                when x"1B6" => data <= "00011";
                when x"1B7" => data <= "00000";
                when x"1B8" => data <= "00000";
                when x"1B9" => data <= "00111";
                when x"1BA" => data <= "01101";
                when x"1BB" => data <= "00110";
                when x"1BC" => data <= "01111";
                when x"1BD" => data <= "01101";
                when x"1BE" => data <= "00000";
                when x"1BF" => data <= "10110";
                when x"1C0" => data <= "00110";
                when x"1C1" => data <= "00000";
                when x"1C2" => data <= "00000";
                when x"1C3" => data <= "00110";
                when x"1C4" => data <= "10110";
                when x"1C5" => data <= "00110";
                when x"1C6" => data <= "00110";
                when x"1C7" => data <= "00110";
                when x"1C8" => data <= "00000";
                when x"1C9" => data <= "00110";
                when x"1CA" => data <= "00000";
                when x"1CB" => data <= "00000";
                when x"1CC" => data <= "00110";
                when x"1CD" => data <= "00000";
                when x"1CE" => data <= "00000";
                when x"1CF" => data <= "00000";
                when x"1D0" => data <= "00110";
                when x"1D1" => data <= "00000";
                when x"1D2" => data <= "00001";
                when x"1D3" => data <= "00000";
                when x"1D4" => data <= "01011";
                when x"1D5" => data <= "00000";
                when x"1D6" => data <= "00000";
                when x"1D7" => data <= "00000";
                when x"1D8" => data <= "00110";
                when x"1D9" => data <= "00111";
                when x"1DA" => data <= "00000";
                when x"1DB" => data <= "00110";
                when x"1DC" => data <= "00110";
                when x"1DD" => data <= "00000";
                when x"1DE" => data <= "00000";
                when x"1DF" => data <= "00110";
                when x"1E0" => data <= "11110";
                when x"1E1" => data <= "00001";
                when x"1E2" => data <= "00110";
                when x"1E3" => data <= "01011";
                when x"1E4" => data <= "00110";
                when x"1E5" => data <= "00000";
                when x"1E6" => data <= "00000";
                when x"1E7" => data <= "01011";
                when x"1E8" => data <= "00000";
                when x"1E9" => data <= "00000";
                when x"1EA" => data <= "00110";
                when x"1EB" => data <= "00110";
                when x"1EC" => data <= "00000";
                when x"1ED" => data <= "10011";
                when x"1EE" => data <= "00110";
                when x"1EF" => data <= "00000";
                when x"1F0" => data <= "00110";
                when x"1F1" => data <= "00110";
                when x"1F2" => data <= "00110";
                when x"1F3" => data <= "00110";
                when x"1F4" => data <= "00000";
                when x"1F5" => data <= "00110";
                when x"1F6" => data <= "10001";
                when x"1F7" => data <= "00110";
                when x"1F8" => data <= "00000";
                when x"1F9" => data <= "00000";
                when x"1FA" => data <= "00110";
                when x"1FB" => data <= "00000";
                when x"1FC" => data <= "00110";
                when x"1FD" => data <= "00000";
                when x"1FE" => data <= "00000";
                when x"1FF" => data <= "00000";
                when x"200" => data <= "00110";
                when x"201" => data <= "00000";
                when x"202" => data <= "11110";
                when x"203" => data <= "00110";
                when x"204" => data <= "00000";
                when x"205" => data <= "00110";
                when x"206" => data <= "00110";
                when x"207" => data <= "00110";
                when x"208" => data <= "00000";
                when x"209" => data <= "00000";
                when x"20A" => data <= "00000";
                when x"20B" => data <= "00110";
                when x"20C" => data <= "01100";
                when x"20D" => data <= "00110";
                when x"20E" => data <= "00110";
                when x"20F" => data <= "00110";
                when x"210" => data <= "11011";
                when x"211" => data <= "00110";
                when x"212" => data <= "00110";
                when x"213" => data <= "00110";
                when x"214" => data <= "00110";
                when x"215" => data <= "00000";
                when x"216" => data <= "11011";
                when x"217" => data <= "10101";
                when x"218" => data <= "00110";
                when x"219" => data <= "00000";
                when x"21A" => data <= "00000";
                when x"21B" => data <= "00000";
                when x"21C" => data <= "00110";
                when x"21D" => data <= "11100";
                when x"21E" => data <= "00000";
                when x"21F" => data <= "00110";
                when x"220" => data <= "00000";
                when x"221" => data <= "00000";
                when x"222" => data <= "00000";
                when x"223" => data <= "00000";
                when x"224" => data <= "00000";
                when x"225" => data <= "00000";
                when x"226" => data <= "00110";
                when x"227" => data <= "00000";
                when x"228" => data <= "00110";
                when x"229" => data <= "00000";
                when x"22A" => data <= "00000";
                when x"22B" => data <= "00000";
                when x"22C" => data <= "10010";
                when x"22D" => data <= "00110";
                when x"22E" => data <= "00100";
                when x"22F" => data <= "00000";
                when x"230" => data <= "00000";
                when x"231" => data <= "00110";
                when x"232" => data <= "01000";
                when x"233" => data <= "00000";
                when x"234" => data <= "00110";
                when x"235" => data <= "00110";
                when x"236" => data <= "01000";
                when x"237" => data <= "01011";
                when x"238" => data <= "10001";
                when x"239" => data <= "00101";
                when x"23A" => data <= "00000";
                when x"23B" => data <= "00000";
                when x"23C" => data <= "00000";
                when x"23D" => data <= "00110";
                when x"23E" => data <= "00000";
                when x"23F" => data <= "00110";
                when x"240" => data <= "00000";
                when x"241" => data <= "00000";
                when x"242" => data <= "00000";
                when x"243" => data <= "00000";
                when x"244" => data <= "00000";
                when x"245" => data <= "00110";
                when x"246" => data <= "00000";
                when x"247" => data <= "00000";
                when x"248" => data <= "00110";
                when x"249" => data <= "00000";
                when x"24A" => data <= "00000";
                when x"24B" => data <= "00110";
                when x"24C" => data <= "00000";
                when x"24D" => data <= "00000";
                when x"24E" => data <= "00000";
                when x"24F" => data <= "01011";
                when x"250" => data <= "00110";
                when x"251" => data <= "11001";
                when x"252" => data <= "11010";
                when x"253" => data <= "00000";
                when x"254" => data <= "00000";
                when x"255" => data <= "00110";
                when x"256" => data <= "00000";
                when x"257" => data <= "00000";
                when x"258" => data <= "00111";
                when x"259" => data <= "00000";
                when x"25A" => data <= "11000";
                when x"25B" => data <= "11010";
                when x"25C" => data <= "00011";
                when x"25D" => data <= "00000";
                when x"25E" => data <= "00000";
                when x"25F" => data <= "00000";
                when x"260" => data <= "00000";
                when x"261" => data <= "01110";
                when x"262" => data <= "00110";
                when x"263" => data <= "00110";
                when x"264" => data <= "00000";
                when x"265" => data <= "11000";
                when x"266" => data <= "00000";
                when x"267" => data <= "00000";
                when x"268" => data <= "00110";
                when x"269" => data <= "00110";
                when x"26A" => data <= "00110";
                when x"26B" => data <= "00000";
                when x"26C" => data <= "10100";
                when x"26D" => data <= "00000";
                when x"26E" => data <= "00100";
                when x"26F" => data <= "01111";
                when x"270" => data <= "00000";
                when x"271" => data <= "00110";
                when x"272" => data <= "00000";
                when x"273" => data <= "00110";
                when x"274" => data <= "00110";
                when x"275" => data <= "00000";
                when x"276" => data <= "11110";
                when x"277" => data <= "00000";
                when x"278" => data <= "00000";
                when x"279" => data <= "00000";
                when x"27A" => data <= "00110";
                when x"27B" => data <= "00110";
                when x"27C" => data <= "00000";
                when x"27D" => data <= "00000";
                when x"27E" => data <= "00110";
                when x"27F" => data <= "10011";
                when x"280" => data <= "00110";
                when x"281" => data <= "00110";
                when x"282" => data <= "11110";
                when x"283" => data <= "00000";
                when x"284" => data <= "00110";
                when x"285" => data <= "00110";
                when x"286" => data <= "00110";
                when x"287" => data <= "00000";
                when x"288" => data <= "00000";
                when x"289" => data <= "00000";
                when x"28A" => data <= "00110";
                when x"28B" => data <= "00110";
                when x"28C" => data <= "00110";
                when x"28D" => data <= "00000";
                when x"28E" => data <= "00100";
                when x"28F" => data <= "00110";
                when x"290" => data <= "11100";
                when x"291" => data <= "01010";
                when x"292" => data <= "00000";
                when x"293" => data <= "00000";
                when x"294" => data <= "00000";
                when x"295" => data <= "00000";
                when x"296" => data <= "00010";
                when x"297" => data <= "00100";
                when x"298" => data <= "00110";
                when x"299" => data <= "00110";
                when x"29A" => data <= "00110";
                when x"29B" => data <= "00110";
                when x"29C" => data <= "00000";
                when x"29D" => data <= "01000";
                when x"29E" => data <= "00000";
                when x"29F" => data <= "10110";
                when x"2A0" => data <= "00000";
                when x"2A1" => data <= "00000";
                when x"2A2" => data <= "00000";
                when x"2A3" => data <= "00110";
                when x"2A4" => data <= "01100";
                when x"2A5" => data <= "11001";
                when x"2A6" => data <= "10001";
                when x"2A7" => data <= "00000";
                when x"2A8" => data <= "00110";
                when x"2A9" => data <= "00000";
                when x"2AA" => data <= "00000";
                when x"2AB" => data <= "11110";
                when x"2AC" => data <= "00110";
                when x"2AD" => data <= "00000";
                when x"2AE" => data <= "00110";
                when x"2AF" => data <= "00000";
                when x"2B0" => data <= "00110";
                when x"2B1" => data <= "00110";
                when x"2B2" => data <= "00110";
                when x"2B3" => data <= "00110";
                when x"2B4" => data <= "00000";
                when x"2B5" => data <= "00110";
                when x"2B6" => data <= "00000";
                when x"2B7" => data <= "00000";
                when x"2B8" => data <= "00110";
                when x"2B9" => data <= "00000";
                when x"2BA" => data <= "00000";
                when x"2BB" => data <= "00000";
                when x"2BC" => data <= "00000";
                when x"2BD" => data <= "00110";
                when x"2BE" => data <= "01101";
                when x"2BF" => data <= "00110";
                when x"2C0" => data <= "00110";
                when x"2C1" => data <= "00110";
                when x"2C2" => data <= "01101";
                when x"2C3" => data <= "00110";
                when x"2C4" => data <= "00000";
                when x"2C5" => data <= "00110";
                when x"2C6" => data <= "00110";
                when x"2C7" => data <= "00000";
                when x"2C8" => data <= "00110";
                when x"2C9" => data <= "00000";
                when x"2CA" => data <= "00000";
                when x"2CB" => data <= "00000";
                when x"2CC" => data <= "00001";
                when x"2CD" => data <= "00110";
                when x"2CE" => data <= "00110";
                when x"2CF" => data <= "01000";
                when x"2D0" => data <= "00110";
                when x"2D1" => data <= "00110";
                when x"2D2" => data <= "00000";
                when x"2D3" => data <= "00110";
                when x"2D4" => data <= "00110";
                when x"2D5" => data <= "00000";
                when x"2D6" => data <= "00000";
                when x"2D7" => data <= "00000";
                when x"2D8" => data <= "00000";
                when x"2D9" => data <= "00110";
                when x"2DA" => data <= "00110";
                when x"2DB" => data <= "00110";
                when x"2DC" => data <= "01011";
                when x"2DD" => data <= "00110";
                when x"2DE" => data <= "00000";
                when x"2DF" => data <= "00000";
                when x"2E0" => data <= "10011";
                when x"2E1" => data <= "10011";
                when x"2E2" => data <= "00000";
                when x"2E3" => data <= "00000";
                when x"2E4" => data <= "00110";
                when x"2E5" => data <= "00000";
                when x"2E6" => data <= "00110";
                when x"2E7" => data <= "00000";
                when x"2E8" => data <= "11001";
                when x"2E9" => data <= "00110";
                when x"2EA" => data <= "00110";
                when x"2EB" => data <= "00100";
                when x"2EC" => data <= "10101";
                when x"2ED" => data <= "00000";
                when x"2EE" => data <= "00110";
                when x"2EF" => data <= "00110";
                when x"2F0" => data <= "00000";
                when x"2F1" => data <= "00000";
                when x"2F2" => data <= "00000";
                when x"2F3" => data <= "11010";
                when x"2F4" => data <= "00110";
                when x"2F5" => data <= "00000";
                when x"2F6" => data <= "00000";
                when x"2F7" => data <= "00000";
                when x"2F8" => data <= "00000";
                when x"2F9" => data <= "00000";
                when x"2FA" => data <= "00000";
                when x"2FB" => data <= "00000";
                when x"2FC" => data <= "01010";
                when x"2FD" => data <= "00110";
                when x"2FE" => data <= "00110";
                when x"2FF" => data <= "00110";
                when x"300" => data <= "00000";
                when x"301" => data <= "01101";
                when x"302" => data <= "00000";
                when x"303" => data <= "11111";
                when x"304" => data <= "00001";
                when x"305" => data <= "11001";
                when x"306" => data <= "00001";
                when x"307" => data <= "00110";
                when x"308" => data <= "11011";
                when x"309" => data <= "00110";
                when x"30A" => data <= "00000";
                when x"30B" => data <= "00110";
                when x"30C" => data <= "00110";
                when x"30D" => data <= "10101";
                when x"30E" => data <= "00000";
                when x"30F" => data <= "11101";
                when x"310" => data <= "00000";
                when x"311" => data <= "00000";
                when x"312" => data <= "00000";
                when x"313" => data <= "00110";
                when x"314" => data <= "01011";
                when x"315" => data <= "00000";
                when x"316" => data <= "00110";
                when x"317" => data <= "11110";
                when x"318" => data <= "00110";
                when x"319" => data <= "00110";
                when x"31A" => data <= "00110";
                when x"31B" => data <= "00110";
                when x"31C" => data <= "00110";
                when x"31D" => data <= "00000";
                when x"31E" => data <= "00000";
                when x"31F" => data <= "00000";
                when x"320" => data <= "00110";
                when x"321" => data <= "00000";
                when x"322" => data <= "00110";
                when x"323" => data <= "00000";
                when x"324" => data <= "00000";
                when x"325" => data <= "00000";
                when x"326" => data <= "11111";
                when x"327" => data <= "00110";
                when x"328" => data <= "00000";
                when x"329" => data <= "00110";
                when x"32A" => data <= "11111";
                when x"32B" => data <= "00110";
                when x"32C" => data <= "00110";
                when x"32D" => data <= "00110";
                when x"32E" => data <= "00000";
                when x"32F" => data <= "10101";
                when x"330" => data <= "00110";
                when x"331" => data <= "00000";
                when x"332" => data <= "00000";
                when x"333" => data <= "00110";
                when x"334" => data <= "00000";
                when x"335" => data <= "00000";
                when x"336" => data <= "00110";
                when x"337" => data <= "11111";
                when x"338" => data <= "00110";
                when x"339" => data <= "00000";
                when x"33A" => data <= "00110";
                when x"33B" => data <= "00110";
                when x"33C" => data <= "00110";
                when x"33D" => data <= "00000";
                when x"33E" => data <= "01011";
                when x"33F" => data <= "00000";
                when x"340" => data <= "00110";
                when x"341" => data <= "00110";
                when x"342" => data <= "00110";
                when x"343" => data <= "00000";
                when x"344" => data <= "00000";
                when x"345" => data <= "11001";
                when x"346" => data <= "10001";
                when x"347" => data <= "00000";
                when x"348" => data <= "00000";
                when x"349" => data <= "10101";
                when x"34A" => data <= "00000";
                when x"34B" => data <= "00000";
                when x"34C" => data <= "00110";
                when x"34D" => data <= "00000";
                when x"34E" => data <= "00110";
                when x"34F" => data <= "00110";
                when x"350" => data <= "11111";
                when x"351" => data <= "00000";
                when x"352" => data <= "00110";
                when x"353" => data <= "00110";
                when x"354" => data <= "00110";
                when x"355" => data <= "01110";
                when x"356" => data <= "00100";
                when x"357" => data <= "00110";
                when x"358" => data <= "00110";
                when x"359" => data <= "00110";
                when x"35A" => data <= "00000";
                when x"35B" => data <= "00110";
                when x"35C" => data <= "00110";
                when x"35D" => data <= "00110";
                when x"35E" => data <= "01101";
                when x"35F" => data <= "00000";
                when x"360" => data <= "00000";
                when x"361" => data <= "00000";
                when x"362" => data <= "01011";
                when x"363" => data <= "00110";
                when x"364" => data <= "00000";
                when x"365" => data <= "00110";
                when x"366" => data <= "01111";
                when x"367" => data <= "00110";
                when x"368" => data <= "00000";
                when x"369" => data <= "00101";
                when x"36A" => data <= "00000";
                when x"36B" => data <= "00110";
                when x"36C" => data <= "00000";
                when x"36D" => data <= "00110";
                when x"36E" => data <= "00000";
                when x"36F" => data <= "01101";
                when x"370" => data <= "00110";
                when x"371" => data <= "10111";
                when x"372" => data <= "00000";
                when x"373" => data <= "00110";
                when x"374" => data <= "00000";
                when x"375" => data <= "00000";
                when x"376" => data <= "00000";
                when x"377" => data <= "00110";
                when x"378" => data <= "00000";
                when x"379" => data <= "01111";
                when x"37A" => data <= "00110";
                when x"37B" => data <= "00110";
                when x"37C" => data <= "00110";
                when x"37D" => data <= "01101";
                when x"37E" => data <= "00000";
                when x"37F" => data <= "01100";
                when x"380" => data <= "00110";
                when x"381" => data <= "00000";
                when x"382" => data <= "00000";
                when x"383" => data <= "00000";
                when x"384" => data <= "00000";
                when x"385" => data <= "00110";
                when x"386" => data <= "00110";
                when x"387" => data <= "00110";
                when x"388" => data <= "00110";
                when x"389" => data <= "00110";
                when x"38A" => data <= "00110";
                when x"38B" => data <= "00110";
                when x"38C" => data <= "00110";
                when x"38D" => data <= "00110";
                when x"38E" => data <= "10101";
                when x"38F" => data <= "00110";
                when x"390" => data <= "00110";
                when x"391" => data <= "10101";
                when x"392" => data <= "01100";
                when x"393" => data <= "00110";
                when x"394" => data <= "01011";
                when x"395" => data <= "00110";
                when x"396" => data <= "00100";
                when x"397" => data <= "01011";
                when x"398" => data <= "00000";
                when x"399" => data <= "00000";
                when x"39A" => data <= "00110";
                when x"39B" => data <= "10010";
                when x"39C" => data <= "00000";
                when x"39D" => data <= "00000";
                when x"39E" => data <= "00000";
                when x"39F" => data <= "00000";
                when x"3A0" => data <= "00000";
                when x"3A1" => data <= "00000";
                when x"3A2" => data <= "00000";
                when x"3A3" => data <= "01011";
                when x"3A4" => data <= "01110";
                when x"3A5" => data <= "00110";
                when x"3A6" => data <= "00101";
                when x"3A7" => data <= "00000";
                when x"3A8" => data <= "10101";
                when x"3A9" => data <= "00110";
                when x"3AA" => data <= "11001";
                when x"3AB" => data <= "00000";
                when x"3AC" => data <= "10101";
                when x"3AD" => data <= "00110";
                when x"3AE" => data <= "00000";
                when x"3AF" => data <= "00000";
                when x"3B0" => data <= "00110";
                when x"3B1" => data <= "00110";
                when x"3B2" => data <= "10010";
                when x"3B3" => data <= "00110";
                when x"3B4" => data <= "00000";
                when x"3B5" => data <= "00000";
                when x"3B6" => data <= "00000";
                when x"3B7" => data <= "00110";
                when x"3B8" => data <= "00011";
                when x"3B9" => data <= "00000";
                when x"3BA" => data <= "00110";
                when x"3BB" => data <= "00110";
                when x"3BC" => data <= "00110";
                when x"3BD" => data <= "00110";
                when x"3BE" => data <= "00110";
                when x"3BF" => data <= "00110";
                when x"3C0" => data <= "01001";
                when x"3C1" => data <= "11001";
                when x"3C2" => data <= "00110";
                when x"3C3" => data <= "10101";
                when x"3C4" => data <= "00000";
                when x"3C5" => data <= "00000";
                when x"3C6" => data <= "00000";
                when x"3C7" => data <= "00000";
                when x"3C8" => data <= "00000";
                when x"3C9" => data <= "00111";
                when x"3CA" => data <= "00000";
                when x"3CB" => data <= "00000";
                when x"3CC" => data <= "10101";
                when x"3CD" => data <= "00000";
                when x"3CE" => data <= "00110";
                when x"3CF" => data <= "01100";
                when x"3D0" => data <= "00110";
                when x"3D1" => data <= "00000";
                when x"3D2" => data <= "00110";
                when x"3D3" => data <= "01001";
                when x"3D4" => data <= "00000";
                when x"3D5" => data <= "00110";
                when x"3D6" => data <= "00000";
                when x"3D7" => data <= "01100";
                when x"3D8" => data <= "00000";
                when x"3D9" => data <= "00000";
                when x"3DA" => data <= "00000";
                when x"3DB" => data <= "00110";
                when x"3DC" => data <= "00110";
                when x"3DD" => data <= "00000";
                when x"3DE" => data <= "00110";
                when x"3DF" => data <= "00001";
                when x"3E0" => data <= "00110";
                when x"3E1" => data <= "00000";
                when x"3E2" => data <= "01111";
                when x"3E3" => data <= "00110";
                when x"3E4" => data <= "00000";
                when x"3E5" => data <= "10011";
                when x"3E6" => data <= "00110";
                when x"3E7" => data <= "00010";
                when x"3E8" => data <= "00110";
                when x"3E9" => data <= "00000";
                when x"3EA" => data <= "00000";
                when x"3EB" => data <= "00110";
                when x"3EC" => data <= "00000";
                when x"3ED" => data <= "00000";
                when x"3EE" => data <= "00110";
                when x"3EF" => data <= "10000";
                when x"3F0" => data <= "00000";
                when x"3F1" => data <= "00111";
                when x"3F2" => data <= "11110";
                when x"3F3" => data <= "00110";
                when x"3F4" => data <= "00110";
                when x"3F5" => data <= "01101";
                when x"3F6" => data <= "00000";
                when x"3F7" => data <= "00000";
                when x"3F8" => data <= "00000";
                when x"3F9" => data <= "00000";
                when x"3FA" => data <= "11111";
                when x"3FB" => data <= "00000";
                when x"3FC" => data <= "00110";
                when x"3FD" => data <= "11011";
                when x"3FE" => data <= "00110";
                when x"3FF" => data <= "11000";
                when x"400" => data <= "00000";
                when x"401" => data <= "00100";
                when x"402" => data <= "00110";
                when x"403" => data <= "00000";
                when x"404" => data <= "10100";
                when x"405" => data <= "00000";
                when x"406" => data <= "00110";
                when x"407" => data <= "01011";
                when x"408" => data <= "00000";
                when x"409" => data <= "00000";
                when x"40A" => data <= "00110";
                when x"40B" => data <= "00110";
                when x"40C" => data <= "00000";
                when x"40D" => data <= "00000";
                when x"40E" => data <= "10000";
                when x"40F" => data <= "00110";
                when x"410" => data <= "10111";
                when x"411" => data <= "00000";
                when x"412" => data <= "01010";
                when x"413" => data <= "00000";
                when x"414" => data <= "00110";
                when x"415" => data <= "00000";
                when x"416" => data <= "00110";
                when x"417" => data <= "11001";
                when x"418" => data <= "01001";
                when x"419" => data <= "00110";
                when x"41A" => data <= "11101";
                when x"41B" => data <= "00000";
                when x"41C" => data <= "10111";
                when x"41D" => data <= "11001";
                when x"41E" => data <= "00000";
                when x"41F" => data <= "00000";
                when x"420" => data <= "10001";
                when x"421" => data <= "00000";
                when x"422" => data <= "11001";
                when x"423" => data <= "00000";
                when x"424" => data <= "10001";
                when x"425" => data <= "00000";
                when x"426" => data <= "10110";
                when x"427" => data <= "00000";
                when x"428" => data <= "00000";
                when x"429" => data <= "00000";
                when x"42A" => data <= "00001";
                when x"42B" => data <= "00000";
                when x"42C" => data <= "10001";
                when x"42D" => data <= "00110";
                when x"42E" => data <= "00000";
                when x"42F" => data <= "00000";
                when x"430" => data <= "00110";
                when x"431" => data <= "00110";
                when x"432" => data <= "00000";
                when x"433" => data <= "00000";
                when x"434" => data <= "00110";
                when x"435" => data <= "00110";
                when x"436" => data <= "11100";
                when x"437" => data <= "00000";
                when x"438" => data <= "00000";
                when x"439" => data <= "00000";
                when x"43A" => data <= "00110";
                when x"43B" => data <= "00000";
                when x"43C" => data <= "00000";
                when x"43D" => data <= "00010";
                when x"43E" => data <= "00000";
                when x"43F" => data <= "10101";
                when x"440" => data <= "00000";
                when x"441" => data <= "00000";
                when x"442" => data <= "00110";
                when x"443" => data <= "00110";
                when x"444" => data <= "00110";
                when x"445" => data <= "01011";
                when x"446" => data <= "11100";
                when x"447" => data <= "00000";
                when x"448" => data <= "00000";
                when x"449" => data <= "00110";
                when x"44A" => data <= "00110";
                when x"44B" => data <= "00000";
                when x"44C" => data <= "00000";
                when x"44D" => data <= "00110";
                when x"44E" => data <= "00000";
                when x"44F" => data <= "00000";
                when x"450" => data <= "00110";
                when x"451" => data <= "01011";
                when x"452" => data <= "00110";
                when x"453" => data <= "00100";
                when x"454" => data <= "00000";
                when x"455" => data <= "00000";
                when x"456" => data <= "01101";
                when x"457" => data <= "00000";
                when x"458" => data <= "00000";
                when x"459" => data <= "11001";
                when x"45A" => data <= "11001";
                when x"45B" => data <= "00110";
                when x"45C" => data <= "00000";
                when x"45D" => data <= "00110";
                when x"45E" => data <= "00110";
                when x"45F" => data <= "00000";
                when x"460" => data <= "00000";
                when x"461" => data <= "00000";
                when x"462" => data <= "00000";
                when x"463" => data <= "00111";
                when x"464" => data <= "00110";
                when x"465" => data <= "00110";
                when x"466" => data <= "10010";
                when x"467" => data <= "00110";
                when x"468" => data <= "01000";
                when x"469" => data <= "00110";
                when x"46A" => data <= "00110";
                when x"46B" => data <= "00110";
                when x"46C" => data <= "00010";
                when x"46D" => data <= "00011";
                when x"46E" => data <= "00110";
                when x"46F" => data <= "00110";
                when x"470" => data <= "00110";
                when x"471" => data <= "00110";
                when x"472" => data <= "00110";
                when x"473" => data <= "00110";
                when x"474" => data <= "00000";
                when x"475" => data <= "00000";
                when x"476" => data <= "00110";
                when x"477" => data <= "11111";
                when x"478" => data <= "00110";
                when x"479" => data <= "10110";
                when x"47A" => data <= "00110";
                when x"47B" => data <= "00110";
                when x"47C" => data <= "00000";
                when x"47D" => data <= "00000";
                when x"47E" => data <= "00110";
                when x"47F" => data <= "00110";
                when x"480" => data <= "00000";
                when x"481" => data <= "00110";
                when x"482" => data <= "00110";
                when x"483" => data <= "00110";
                when x"484" => data <= "00110";
                when x"485" => data <= "00110";
                when x"486" => data <= "01101";
                when x"487" => data <= "01000";
                when x"488" => data <= "00110";
                when x"489" => data <= "00000";
                when x"48A" => data <= "01111";
                when x"48B" => data <= "10011";
                when x"48C" => data <= "10111";
                when x"48D" => data <= "00110";
                when x"48E" => data <= "00110";
                when x"48F" => data <= "00110";
                when x"490" => data <= "00000";
                when x"491" => data <= "01011";
                when x"492" => data <= "00110";
                when x"493" => data <= "00000";
                when x"494" => data <= "00000";
                when x"495" => data <= "00000";
                when x"496" => data <= "00000";
                when x"497" => data <= "00110";
                when x"498" => data <= "00000";
                when x"499" => data <= "11010";
                when x"49A" => data <= "00000";
                when x"49B" => data <= "00110";
                when x"49C" => data <= "00000";
                when x"49D" => data <= "11100";
                when x"49E" => data <= "00110";
                when x"49F" => data <= "00000";
                when x"4A0" => data <= "00110";
                when x"4A1" => data <= "00000";
                when x"4A2" => data <= "00110";
                when x"4A3" => data <= "00000";
                when x"4A4" => data <= "01100";
                when x"4A5" => data <= "11010";
                when x"4A6" => data <= "00000";
                when x"4A7" => data <= "00000";
                when x"4A8" => data <= "00000";
                when x"4A9" => data <= "00000";
                when x"4AA" => data <= "00110";
                when x"4AB" => data <= "00000";
                when x"4AC" => data <= "10111";
                when x"4AD" => data <= "11001";
                when x"4AE" => data <= "00000";
                when x"4AF" => data <= "00000";
                when x"4B0" => data <= "00110";
                when x"4B1" => data <= "00110";
                when x"4B2" => data <= "00110";
                when x"4B3" => data <= "00000";
                when x"4B4" => data <= "00110";
                when x"4B5" => data <= "00100";
                when x"4B6" => data <= "00110";
                when x"4B7" => data <= "00000";
                when x"4B8" => data <= "00000";
                when x"4B9" => data <= "00110";
                when x"4BA" => data <= "00000";
                when x"4BB" => data <= "00000";
                when x"4BC" => data <= "00000";
                when x"4BD" => data <= "00000";
                when x"4BE" => data <= "00110";
                when x"4BF" => data <= "00000";
                when x"4C0" => data <= "00000";
                when x"4C1" => data <= "00000";
                when x"4C2" => data <= "00000";
                when x"4C3" => data <= "00000";
                when x"4C4" => data <= "00000";
                when x"4C5" => data <= "00110";
                when x"4C6" => data <= "00110";
                when x"4C7" => data <= "00000";
                when x"4C8" => data <= "00000";
                when x"4C9" => data <= "00000";
                when x"4CA" => data <= "01101";
                when x"4CB" => data <= "00000";
                when x"4CC" => data <= "00000";
                when x"4CD" => data <= "00000";
                when x"4CE" => data <= "00000";
                when x"4CF" => data <= "00110";
                when x"4D0" => data <= "00000";
                when x"4D1" => data <= "00000";
                when x"4D2" => data <= "00110";
                when x"4D3" => data <= "00110";
                when x"4D4" => data <= "00110";
                when x"4D5" => data <= "00000";
                when x"4D6" => data <= "00110";
                when x"4D7" => data <= "00000";
                when x"4D8" => data <= "01011";
                when x"4D9" => data <= "11110";
                when x"4DA" => data <= "00000";
                when x"4DB" => data <= "00110";
                when x"4DC" => data <= "01011";
                when x"4DD" => data <= "00110";
                when x"4DE" => data <= "00110";
                when x"4DF" => data <= "00000";
                when x"4E0" => data <= "00110";
                when x"4E1" => data <= "10001";
                when x"4E2" => data <= "01100";
                when x"4E3" => data <= "01000";
                when x"4E4" => data <= "00000";
                when x"4E5" => data <= "00110";
                when x"4E6" => data <= "00000";
                when x"4E7" => data <= "00000";
                when x"4E8" => data <= "10010";
                when x"4E9" => data <= "00000";
                when x"4EA" => data <= "00000";
                when x"4EB" => data <= "00110";
                when x"4EC" => data <= "00000";
                when x"4ED" => data <= "10010";
                when x"4EE" => data <= "00000";
                when x"4EF" => data <= "00000";
                when x"4F0" => data <= "00110";
                when x"4F1" => data <= "00110";
                when x"4F2" => data <= "00110";
                when x"4F3" => data <= "00000";
                when x"4F4" => data <= "00110";
                when x"4F5" => data <= "01110";
                when x"4F6" => data <= "00110";
                when x"4F7" => data <= "00000";
                when x"4F8" => data <= "00110";
                when x"4F9" => data <= "00000";
                when x"4FA" => data <= "10010";
                when x"4FB" => data <= "00110";
                when x"4FC" => data <= "00110";
                when x"4FD" => data <= "00000";
                when x"4FE" => data <= "00110";
                when x"4FF" => data <= "00000";
                when x"500" => data <= "00000";
                when x"501" => data <= "11000";
                when x"502" => data <= "00110";
                when x"503" => data <= "00000";
                when x"504" => data <= "00110";
                when x"505" => data <= "00000";
                when x"506" => data <= "01001";
                when x"507" => data <= "00000";
                when x"508" => data <= "00110";
                when x"509" => data <= "00110";
                when x"50A" => data <= "00110";
                when x"50B" => data <= "10010";
                when x"50C" => data <= "00110";
                when x"50D" => data <= "01111";
                when x"50E" => data <= "10011";
                when x"50F" => data <= "01101";
                when x"510" => data <= "00111";
                when x"511" => data <= "01101";
                when x"512" => data <= "00000";
                when x"513" => data <= "00110";
                when x"514" => data <= "00110";
                when x"515" => data <= "00110";
                when x"516" => data <= "00000";
                when x"517" => data <= "00110";
                when x"518" => data <= "00000";
                when x"519" => data <= "00000";
                when x"51A" => data <= "00110";
                when x"51B" => data <= "01111";
                when x"51C" => data <= "00000";
                when x"51D" => data <= "00000";
                when x"51E" => data <= "00000";
                when x"51F" => data <= "10100";
                when x"520" => data <= "00110";
                when x"521" => data <= "00000";
                when x"522" => data <= "01000";
                when x"523" => data <= "00110";
                when x"524" => data <= "11111";
                when x"525" => data <= "11001";
                when x"526" => data <= "00110";
                when x"527" => data <= "00110";
                when x"528" => data <= "10101";
                when x"529" => data <= "00110";
                when x"52A" => data <= "00110";
                when x"52B" => data <= "00000";
                when x"52C" => data <= "00110";
                when x"52D" => data <= "00110";
                when x"52E" => data <= "00000";
                when x"52F" => data <= "00000";
                when x"530" => data <= "00000";
                when x"531" => data <= "10100";
                when x"532" => data <= "11100";
                when x"533" => data <= "01011";
                when x"534" => data <= "00000";
                when x"535" => data <= "00000";
                when x"536" => data <= "00110";
                when x"537" => data <= "00110";
                when x"538" => data <= "00110";
                when x"539" => data <= "11010";
                when x"53A" => data <= "00000";
                when x"53B" => data <= "00100";
                when x"53C" => data <= "00110";
                when x"53D" => data <= "10011";
                when x"53E" => data <= "00110";
                when x"53F" => data <= "11111";
                when x"540" => data <= "00000";
                when x"541" => data <= "00000";
                when x"542" => data <= "00110";
                when x"543" => data <= "00000";
                when x"544" => data <= "00110";
                when x"545" => data <= "00000";
                when x"546" => data <= "10000";
                when x"547" => data <= "00110";
                when x"548" => data <= "01101";
                when x"549" => data <= "00110";
                when x"54A" => data <= "00000";
                when x"54B" => data <= "00110";
                when x"54C" => data <= "00110";
                when x"54D" => data <= "00110";
                when x"54E" => data <= "00000";
                when x"54F" => data <= "11001";
                when x"550" => data <= "00000";
                when x"551" => data <= "01000";
                when x"552" => data <= "00000";
                when x"553" => data <= "00000";
                when x"554" => data <= "00000";
                when x"555" => data <= "00000";
                when x"556" => data <= "00000";
                when x"557" => data <= "00110";
                when x"558" => data <= "00110";
                when x"559" => data <= "00000";
                when x"55A" => data <= "10001";
                when x"55B" => data <= "00110";
                when x"55C" => data <= "00000";
                when x"55D" => data <= "00110";
                when x"55E" => data <= "00100";
                when x"55F" => data <= "01010";
                when x"560" => data <= "00110";
                when x"561" => data <= "00110";
                when x"562" => data <= "00000";
                when x"563" => data <= "01110";
                when x"564" => data <= "00110";
                when x"565" => data <= "00000";
                when x"566" => data <= "01100";
                when x"567" => data <= "00110";
                when x"568" => data <= "00000";
                when x"569" => data <= "00000";
                when x"56A" => data <= "00000";
                when x"56B" => data <= "00110";
                when x"56C" => data <= "00110";
                when x"56D" => data <= "00000";
                when x"56E" => data <= "00000";
                when x"56F" => data <= "00110";
                when x"570" => data <= "01011";
                when x"571" => data <= "00110";
                when x"572" => data <= "00110";
                when x"573" => data <= "11001";
                when x"574" => data <= "00110";
                when x"575" => data <= "00110";
                when x"576" => data <= "00110";
                when x"577" => data <= "00000";
                when x"578" => data <= "00110";
                when x"579" => data <= "00000";
                when x"57A" => data <= "01011";
                when x"57B" => data <= "01110";
                when x"57C" => data <= "00110";
                when x"57D" => data <= "00110";
                when x"57E" => data <= "00000";
                when x"57F" => data <= "00000";
                when x"580" => data <= "10001";
                when x"581" => data <= "11000";
                when x"582" => data <= "00110";
                when x"583" => data <= "00110";
                when x"584" => data <= "00000";
                when x"585" => data <= "00110";
                when x"586" => data <= "00000";
                when x"587" => data <= "00000";
                when x"588" => data <= "11000";
                when x"589" => data <= "00110";
                when x"58A" => data <= "10011";
                when x"58B" => data <= "10001";
                when x"58C" => data <= "00110";
                when x"58D" => data <= "00110";
                when x"58E" => data <= "00000";
                when x"58F" => data <= "11001";
                when x"590" => data <= "00000";
                when x"591" => data <= "00000";
                when x"592" => data <= "00000";
                when x"593" => data <= "00110";
                when x"594" => data <= "00000";
                when x"595" => data <= "11000";
                when x"596" => data <= "01011";
                when x"597" => data <= "00000";
                when x"598" => data <= "00001";
                when x"599" => data <= "00110";
                when x"59A" => data <= "00110";
                when x"59B" => data <= "00110";
                when x"59C" => data <= "00100";
                when x"59D" => data <= "00110";
                when x"59E" => data <= "11100";
                when x"59F" => data <= "00000";
                when x"5A0" => data <= "00000";
                when x"5A1" => data <= "01100";
                when x"5A2" => data <= "00110";
                when x"5A3" => data <= "00110";
                when x"5A4" => data <= "01101";
                when x"5A5" => data <= "00000";
                when x"5A6" => data <= "11001";
                when x"5A7" => data <= "00000";
                when x"5A8" => data <= "00110";
                when x"5A9" => data <= "00110";
                when x"5AA" => data <= "00000";
                when x"5AB" => data <= "01011";
                when x"5AC" => data <= "00110";
                when x"5AD" => data <= "00000";
                when x"5AE" => data <= "00110";
                when x"5AF" => data <= "10111";
                when x"5B0" => data <= "00110";
                when x"5B1" => data <= "00000";
                when x"5B2" => data <= "10001";
                when x"5B3" => data <= "00000";
                when x"5B4" => data <= "00000";
                when x"5B5" => data <= "01011";
                when x"5B6" => data <= "01010";
                when x"5B7" => data <= "00110";
                when x"5B8" => data <= "00110";
                when x"5B9" => data <= "01010";
                when x"5BA" => data <= "00000";
                when x"5BB" => data <= "00110";
                when x"5BC" => data <= "00000";
                when x"5BD" => data <= "00000";
                when x"5BE" => data <= "00000";
                when x"5BF" => data <= "00110";
                when x"5C0" => data <= "00110";
                when x"5C1" => data <= "00110";
                when x"5C2" => data <= "01001";
                when x"5C3" => data <= "01100";
                when x"5C4" => data <= "00000";
                when x"5C5" => data <= "00110";
                when x"5C6" => data <= "00000";
                when x"5C7" => data <= "00110";
                when x"5C8" => data <= "00000";
                when x"5C9" => data <= "11010";
                when x"5CA" => data <= "10101";
                when x"5CB" => data <= "00000";
                when x"5CC" => data <= "00110";
                when x"5CD" => data <= "00000";
                when x"5CE" => data <= "00000";
                when x"5CF" => data <= "00000";
                when x"5D0" => data <= "01011";
                when x"5D1" => data <= "00000";
                when x"5D2" => data <= "11111";
                when x"5D3" => data <= "00000";
                when x"5D4" => data <= "01101";
                when x"5D5" => data <= "00110";
                when x"5D6" => data <= "01011";
                when x"5D7" => data <= "00110";
                when x"5D8" => data <= "10100";
                when x"5D9" => data <= "00000";
                when x"5DA" => data <= "00110";
                when x"5DB" => data <= "00000";
                when x"5DC" => data <= "00110";
                when x"5DD" => data <= "00000";
                when x"5DE" => data <= "00110";
                when x"5DF" => data <= "00110";
                when x"5E0" => data <= "00000";
                when x"5E1" => data <= "01010";
                when x"5E2" => data <= "00000";
                when x"5E3" => data <= "00000";
                when x"5E4" => data <= "00000";
                when x"5E5" => data <= "00000";
                when x"5E6" => data <= "00000";
                when x"5E7" => data <= "00000";
                when x"5E8" => data <= "00000";
                when x"5E9" => data <= "00000";
                when x"5EA" => data <= "11110";
                when x"5EB" => data <= "00000";
                when x"5EC" => data <= "10111";
                when x"5ED" => data <= "00000";
                when x"5EE" => data <= "00000";
                when x"5EF" => data <= "00110";
                when x"5F0" => data <= "00110";
                when x"5F1" => data <= "00000";
                when x"5F2" => data <= "11100";
                when x"5F3" => data <= "00110";
                when x"5F4" => data <= "00000";
                when x"5F5" => data <= "00110";
                when x"5F6" => data <= "11001";
                when x"5F7" => data <= "00110";
                when x"5F8" => data <= "00110";
                when x"5F9" => data <= "00101";
                when x"5FA" => data <= "11101";
                when x"5FB" => data <= "00110";
                when x"5FC" => data <= "00000";
                when x"5FD" => data <= "00000";
                when x"5FE" => data <= "01001";
                when x"5FF" => data <= "01110";
                when x"600" => data <= "00000";
                when x"601" => data <= "00000";
                when x"602" => data <= "00000";
                when x"603" => data <= "00110";
                when x"604" => data <= "00110";
                when x"605" => data <= "00000";
                when x"606" => data <= "01101";
                when x"607" => data <= "10110";
                when x"608" => data <= "11111";
                when x"609" => data <= "00000";
                when x"60A" => data <= "00000";
                when x"60B" => data <= "00110";
                when x"60C" => data <= "00000";
                when x"60D" => data <= "00110";
                when x"60E" => data <= "11001";
                when x"60F" => data <= "00000";
                when x"610" => data <= "00110";
                when x"611" => data <= "00000";
                when x"612" => data <= "11001";
                when x"613" => data <= "00000";
                when x"614" => data <= "00110";
                when x"615" => data <= "00000";
                when x"616" => data <= "00101";
                when x"617" => data <= "11111";
                when x"618" => data <= "11111";
                when x"619" => data <= "00000";
                when x"61A" => data <= "01101";
                when x"61B" => data <= "00110";
                when x"61C" => data <= "00110";
                when x"61D" => data <= "01101";
                when x"61E" => data <= "00110";
                when x"61F" => data <= "00000";
                when x"620" => data <= "00110";
                when x"621" => data <= "00000";
                when x"622" => data <= "00110";
                when x"623" => data <= "00000";
                when x"624" => data <= "00000";
                when x"625" => data <= "00110";
                when x"626" => data <= "11000";
                when x"627" => data <= "00000";
                when x"628" => data <= "00110";
                when x"629" => data <= "10110";
                when x"62A" => data <= "00000";
                when x"62B" => data <= "11001";
                when x"62C" => data <= "10101";
                when x"62D" => data <= "00110";
                when x"62E" => data <= "00110";
                when x"62F" => data <= "00110";
                when x"630" => data <= "00000";
                when x"631" => data <= "00110";
                when x"632" => data <= "00000";
                when x"633" => data <= "00000";
                when x"634" => data <= "01011";
                when x"635" => data <= "00000";
                when x"636" => data <= "00000";
                when x"637" => data <= "00110";
                when x"638" => data <= "00000";
                when x"639" => data <= "00000";
                when x"63A" => data <= "00000";
                when x"63B" => data <= "00110";
                when x"63C" => data <= "00000";
                when x"63D" => data <= "11111";
                when x"63E" => data <= "00000";
                when x"63F" => data <= "01000";
                when x"640" => data <= "00000";
                when x"641" => data <= "01001";
                when x"642" => data <= "00110";
                when x"643" => data <= "00000";
                when x"644" => data <= "00000";
                when x"645" => data <= "00110";
                when x"646" => data <= "00000";
                when x"647" => data <= "11000";
                when x"648" => data <= "00000";
                when x"649" => data <= "00110";
                when x"64A" => data <= "01100";
                when x"64B" => data <= "00000";
                when x"64C" => data <= "00110";
                when x"64D" => data <= "00000";
                when x"64E" => data <= "00000";
                when x"64F" => data <= "11011";
                when x"650" => data <= "00101";
                when x"651" => data <= "00110";
                when x"652" => data <= "00110";
                when x"653" => data <= "00110";
                when x"654" => data <= "00000";
                when x"655" => data <= "00110";
                when x"656" => data <= "00000";
                when x"657" => data <= "00110";
                when x"658" => data <= "00000";
                when x"659" => data <= "01100";
                when x"65A" => data <= "00000";
                when x"65B" => data <= "00110";
                when x"65C" => data <= "00000";
                when x"65D" => data <= "00001";
                when x"65E" => data <= "00110";
                when x"65F" => data <= "00110";
                when x"660" => data <= "00110";
                when x"661" => data <= "00110";
                when x"662" => data <= "00000";
                when x"663" => data <= "00110";
                when x"664" => data <= "01000";
                when x"665" => data <= "00000";
                when x"666" => data <= "00000";
                when x"667" => data <= "01001";
                when x"668" => data <= "00000";
                when x"669" => data <= "00000";
                when x"66A" => data <= "00110";
                when x"66B" => data <= "00000";
                when x"66C" => data <= "00110";
                when x"66D" => data <= "00000";
                when x"66E" => data <= "00000";
                when x"66F" => data <= "11001";
                when x"670" => data <= "00110";
                when x"671" => data <= "11111";
                when x"672" => data <= "00110";
                when x"673" => data <= "00000";
                when x"674" => data <= "00110";
                when x"675" => data <= "00110";
                when x"676" => data <= "00110";
                when x"677" => data <= "11001";
                when x"678" => data <= "00110";
                when x"679" => data <= "00110";
                when x"67A" => data <= "01101";
                when x"67B" => data <= "00000";
                when x"67C" => data <= "00000";
                when x"67D" => data <= "00110";
                when x"67E" => data <= "00110";
                when x"67F" => data <= "00110";
                when x"680" => data <= "00000";
                when x"681" => data <= "00110";
                when x"682" => data <= "00101";
                when x"683" => data <= "00000";
                when x"684" => data <= "00000";
                when x"685" => data <= "00110";
                when x"686" => data <= "00000";
                when x"687" => data <= "00000";
                when x"688" => data <= "00110";
                when x"689" => data <= "00110";
                when x"68A" => data <= "00000";
                when x"68B" => data <= "00000";
                when x"68C" => data <= "00000";
                when x"68D" => data <= "00110";
                when x"68E" => data <= "00000";
                when x"68F" => data <= "00110";
                when x"690" => data <= "00110";
                when x"691" => data <= "00000";
                when x"692" => data <= "00000";
                when x"693" => data <= "00110";
                when x"694" => data <= "00000";
                when x"695" => data <= "00000";
                when x"696" => data <= "00000";
                when x"697" => data <= "00000";
                when x"698" => data <= "00000";
                when x"699" => data <= "00000";
                when x"69A" => data <= "00110";
                when x"69B" => data <= "01111";
                when x"69C" => data <= "00110";
                when x"69D" => data <= "00110";
                when x"69E" => data <= "00010";
                when x"69F" => data <= "00000";
                when x"6A0" => data <= "00110";
                when x"6A1" => data <= "00011";
                when x"6A2" => data <= "00110";
                when x"6A3" => data <= "00000";
                when x"6A4" => data <= "00000";
                when x"6A5" => data <= "00000";
                when x"6A6" => data <= "00110";
                when x"6A7" => data <= "00000";
                when x"6A8" => data <= "00110";
                when x"6A9" => data <= "00000";
                when x"6AA" => data <= "00110";
                when x"6AB" => data <= "00110";
                when x"6AC" => data <= "00110";
                when x"6AD" => data <= "00110";
                when x"6AE" => data <= "01101";
                when x"6AF" => data <= "00000";
                when x"6B0" => data <= "00000";
                when x"6B1" => data <= "00000";
                when x"6B2" => data <= "11101";
                when x"6B3" => data <= "00110";
                when x"6B4" => data <= "00110";
                when x"6B5" => data <= "00000";
                when x"6B6" => data <= "00110";
                when x"6B7" => data <= "00000";
                when x"6B8" => data <= "00000";
                when x"6B9" => data <= "00000";
                when x"6BA" => data <= "00110";
                when x"6BB" => data <= "00000";
                when x"6BC" => data <= "00110";
                when x"6BD" => data <= "00000";
                when x"6BE" => data <= "00000";
                when x"6BF" => data <= "00000";
                when x"6C0" => data <= "00000";
                when x"6C1" => data <= "00000";
                when x"6C2" => data <= "00000";
                when x"6C3" => data <= "00000";
                when x"6C4" => data <= "00110";
                when x"6C5" => data <= "00110";
                when x"6C6" => data <= "00001";
                when x"6C7" => data <= "00110";
                when x"6C8" => data <= "00110";
                when x"6C9" => data <= "00000";
                when x"6CA" => data <= "00110";
                when x"6CB" => data <= "00110";
                when x"6CC" => data <= "11110";
                when x"6CD" => data <= "00000";
                when x"6CE" => data <= "00000";
                when x"6CF" => data <= "00000";
                when x"6D0" => data <= "00000";
                when x"6D1" => data <= "00110";
                when x"6D2" => data <= "00110";
                when x"6D3" => data <= "00000";
                when x"6D4" => data <= "00000";
                when x"6D5" => data <= "00110";
                when x"6D6" => data <= "01001";
                when x"6D7" => data <= "00110";
                when x"6D8" => data <= "00110";
                when x"6D9" => data <= "00110";
                when x"6DA" => data <= "00000";
                when x"6DB" => data <= "00110";
                when x"6DC" => data <= "00110";
                when x"6DD" => data <= "01011";
                when x"6DE" => data <= "00110";
                when x"6DF" => data <= "00110";
                when x"6E0" => data <= "00110";
                when x"6E1" => data <= "00110";
                when x"6E2" => data <= "00000";
                when x"6E3" => data <= "00000";
                when x"6E4" => data <= "00000";
                when x"6E5" => data <= "00110";
                when x"6E6" => data <= "00000";
                when x"6E7" => data <= "00000";
                when x"6E8" => data <= "00000";
                when x"6E9" => data <= "00110";
                when x"6EA" => data <= "00000";
                when x"6EB" => data <= "00110";
                when x"6EC" => data <= "10000";
                when x"6ED" => data <= "00000";
                when x"6EE" => data <= "01101";
                when x"6EF" => data <= "00110";
                when x"6F0" => data <= "00110";
                when x"6F1" => data <= "00000";
                when x"6F2" => data <= "00110";
                when x"6F3" => data <= "00000";
                when x"6F4" => data <= "00000";
                when x"6F5" => data <= "00000";
                when x"6F6" => data <= "00000";
                when x"6F7" => data <= "00000";
                when x"6F8" => data <= "11000";
                when x"6F9" => data <= "00110";
                when x"6FA" => data <= "00000";
                when x"6FB" => data <= "00110";
                when x"6FC" => data <= "00000";
                when x"6FD" => data <= "00000";
                when x"6FE" => data <= "00000";
                when x"6FF" => data <= "00110";
                when x"700" => data <= "00110";
                when x"701" => data <= "00000";
                when x"702" => data <= "00001";
                when x"703" => data <= "00000";
                when x"704" => data <= "00010";
                when x"705" => data <= "10000";
                when x"706" => data <= "00110";
                when x"707" => data <= "00110";
                when x"708" => data <= "00000";
                when x"709" => data <= "00110";
                when x"70A" => data <= "00110";
                when x"70B" => data <= "10111";
                when x"70C" => data <= "00000";
                when x"70D" => data <= "00100";
                when x"70E" => data <= "01100";
                when x"70F" => data <= "11100";
                when x"710" => data <= "00110";
                when x"711" => data <= "00000";
                when x"712" => data <= "01011";
                when x"713" => data <= "11010";
                when x"714" => data <= "00000";
                when x"715" => data <= "01011";
                when x"716" => data <= "00110";
                when x"717" => data <= "01110";
                when x"718" => data <= "00110";
                when x"719" => data <= "10101";
                when x"71A" => data <= "00000";
                when x"71B" => data <= "00110";
                when x"71C" => data <= "00000";
                when x"71D" => data <= "00000";
                when x"71E" => data <= "00110";
                when x"71F" => data <= "00110";
                when x"720" => data <= "00000";
                when x"721" => data <= "11000";
                when x"722" => data <= "01101";
                when x"723" => data <= "00000";
                when x"724" => data <= "00000";
                when x"725" => data <= "11100";
                when x"726" => data <= "00110";
                when x"727" => data <= "00110";
                when x"728" => data <= "00110";
                when x"729" => data <= "00000";
                when x"72A" => data <= "00110";
                when x"72B" => data <= "01101";
                when x"72C" => data <= "00000";
                when x"72D" => data <= "00101";
                when x"72E" => data <= "00110";
                when x"72F" => data <= "00000";
                when x"730" => data <= "00110";
                when x"731" => data <= "00000";
                when x"732" => data <= "00000";
                when x"733" => data <= "10011";
                when x"734" => data <= "00000";
                when x"735" => data <= "00110";
                when x"736" => data <= "00110";
                when x"737" => data <= "00000";
                when x"738" => data <= "00000";
                when x"739" => data <= "00110";
                when x"73A" => data <= "00000";
                when x"73B" => data <= "00110";
                when x"73C" => data <= "10100";
                when x"73D" => data <= "00000";
                when x"73E" => data <= "00000";
                when x"73F" => data <= "00000";
                when x"740" => data <= "00110";
                when x"741" => data <= "00110";
                when x"742" => data <= "00000";
                when x"743" => data <= "00000";
                when x"744" => data <= "00101";
                when x"745" => data <= "00110";
                when x"746" => data <= "00001";
                when x"747" => data <= "00110";
                when x"748" => data <= "01101";
                when x"749" => data <= "00110";
                when x"74A" => data <= "00110";
                when x"74B" => data <= "00001";
                when x"74C" => data <= "00110";
                when x"74D" => data <= "00000";
                when x"74E" => data <= "00110";
                when x"74F" => data <= "00110";
                when x"750" => data <= "00000";
                when x"751" => data <= "00101";
                when x"752" => data <= "00110";
                when x"753" => data <= "00000";
                when x"754" => data <= "00000";
                when x"755" => data <= "10100";
                when x"756" => data <= "00000";
                when x"757" => data <= "00000";
                when x"758" => data <= "00110";
                when x"759" => data <= "00110";
                when x"75A" => data <= "00110";
                when x"75B" => data <= "00000";
                when x"75C" => data <= "01011";
                when x"75D" => data <= "00000";
                when x"75E" => data <= "00000";
                when x"75F" => data <= "00000";
                when x"760" => data <= "00110";
                when x"761" => data <= "11111";
                when x"762" => data <= "00000";
                when x"763" => data <= "00000";
                when x"764" => data <= "00000";
                when x"765" => data <= "00000";
                when x"766" => data <= "00110";
                when x"767" => data <= "00000";
                when x"768" => data <= "00000";
                when x"769" => data <= "00000";
                when x"76A" => data <= "00000";
                when x"76B" => data <= "00000";
                when x"76C" => data <= "00111";
                when x"76D" => data <= "00110";
                when x"76E" => data <= "00000";
                when x"76F" => data <= "00110";
                when x"770" => data <= "00000";
                when x"771" => data <= "00110";
                when x"772" => data <= "00000";
                when x"773" => data <= "10010";
                when x"774" => data <= "00000";
                when x"775" => data <= "00110";
                when x"776" => data <= "11101";
                when x"777" => data <= "00000";
                when x"778" => data <= "00000";
                when x"779" => data <= "00000";
                when x"77A" => data <= "00000";
                when x"77B" => data <= "00000";
                when x"77C" => data <= "00000";
                when x"77D" => data <= "00000";
                when x"77E" => data <= "10011";
                when x"77F" => data <= "00000";
                when x"780" => data <= "00110";
                when x"781" => data <= "01101";
                when x"782" => data <= "00000";
                when x"783" => data <= "00110";
                when x"784" => data <= "00000";
                when x"785" => data <= "00000";
                when x"786" => data <= "00000";
                when x"787" => data <= "00110";
                when x"788" => data <= "01000";
                when x"789" => data <= "00110";
                when x"78A" => data <= "00000";
                when x"78B" => data <= "11001";
                when x"78C" => data <= "00110";
                when x"78D" => data <= "00000";
                when x"78E" => data <= "01010";
                when x"78F" => data <= "01011";
                when x"790" => data <= "11001";
                when x"791" => data <= "00000";
                when x"792" => data <= "00000";
                when x"793" => data <= "00000";
                when x"794" => data <= "00110";
                when x"795" => data <= "10101";
                when x"796" => data <= "00110";
                when x"797" => data <= "00110";
                when x"798" => data <= "00110";
                when x"799" => data <= "00000";
                when x"79A" => data <= "00110";
                when x"79B" => data <= "00000";
                when x"79C" => data <= "00000";
                when x"79D" => data <= "00110";
                when x"79E" => data <= "11100";
                when x"79F" => data <= "00010";
                when x"7A0" => data <= "01101";
                when x"7A1" => data <= "00110";
                when x"7A2" => data <= "00110";
                when x"7A3" => data <= "00000";
                when x"7A4" => data <= "00110";
                when x"7A5" => data <= "00000";
                when x"7A6" => data <= "01001";
                when x"7A7" => data <= "00000";
                when x"7A8" => data <= "00000";
                when x"7A9" => data <= "00000";
                when x"7AA" => data <= "00110";
                when x"7AB" => data <= "00110";
                when x"7AC" => data <= "00000";
                when x"7AD" => data <= "01110";
                when x"7AE" => data <= "00000";
                when x"7AF" => data <= "11010";
                when x"7B0" => data <= "11010";
                when x"7B1" => data <= "00110";
                when x"7B2" => data <= "01011";
                when x"7B3" => data <= "00000";
                when x"7B4" => data <= "00110";
                when x"7B5" => data <= "00110";
                when x"7B6" => data <= "00000";
                when x"7B7" => data <= "00001";
                when x"7B8" => data <= "10111";
                when x"7B9" => data <= "11010";
                when x"7BA" => data <= "00110";
                when x"7BB" => data <= "00000";
                when x"7BC" => data <= "00000";
                when x"7BD" => data <= "11111";
                when x"7BE" => data <= "00000";
                when x"7BF" => data <= "00110";
                when x"7C0" => data <= "00000";
                when x"7C1" => data <= "10010";
                when x"7C2" => data <= "00000";
                when x"7C3" => data <= "00000";
                when x"7C4" => data <= "00110";
                when x"7C5" => data <= "10001";
                when x"7C6" => data <= "00000";
                when x"7C7" => data <= "00110";
                when x"7C8" => data <= "00000";
                when x"7C9" => data <= "01010";
                when x"7CA" => data <= "10110";
                when x"7CB" => data <= "01100";
                when x"7CC" => data <= "00000";
                when x"7CD" => data <= "00110";
                when x"7CE" => data <= "00110";
                when x"7CF" => data <= "10000";
                when x"7D0" => data <= "00000";
                when x"7D1" => data <= "00000";
                when x"7D2" => data <= "00110";
                when x"7D3" => data <= "00110";
                when x"7D4" => data <= "00011";
                when x"7D5" => data <= "01011";
                when x"7D6" => data <= "00000";
                when x"7D7" => data <= "00000";
                when x"7D8" => data <= "01101";
                when x"7D9" => data <= "00110";
                when x"7DA" => data <= "00000";
                when x"7DB" => data <= "01011";
                when x"7DC" => data <= "00000";
                when x"7DD" => data <= "00110";
                when x"7DE" => data <= "00110";
                when x"7DF" => data <= "00110";
                when x"7E0" => data <= "00110";
                when x"7E1" => data <= "00110";
                when x"7E2" => data <= "00000";
                when x"7E3" => data <= "00110";
                when x"7E4" => data <= "00000";
                when x"7E5" => data <= "00000";
                when x"7E6" => data <= "00000";
                when x"7E7" => data <= "00110";
                when x"7E8" => data <= "10101";
                when x"7E9" => data <= "00110";
                when x"7EA" => data <= "00000";
                when x"7EB" => data <= "00110";
                when x"7EC" => data <= "00000";
                when x"7ED" => data <= "00110";
                when x"7EE" => data <= "00110";
                when x"7EF" => data <= "00110";
                when x"7F0" => data <= "00110";
                when x"7F1" => data <= "00110";
                when x"7F2" => data <= "00000";
                when x"7F3" => data <= "00000";
                when x"7F4" => data <= "00000";
                when x"7F5" => data <= "00000";
                when x"7F6" => data <= "00000";
                when x"7F7" => data <= "00000";
                when x"7F8" => data <= "00000";
                when x"7F9" => data <= "00000";
                when x"7FA" => data <= "10001";
                when x"7FB" => data <= "00110";
                when x"7FC" => data <= "11001";
                when x"7FD" => data <= "00110";
                when x"7FE" => data <= "01000";
                when x"7FF" => data <= "00110";
                when x"800" => data <= "00110";
                when x"801" => data <= "00000";
                when x"802" => data <= "00110";
                when x"803" => data <= "00000";
                when x"804" => data <= "00110";
                when x"805" => data <= "00000";
                when x"806" => data <= "00110";
                when x"807" => data <= "00110";
                when x"808" => data <= "00110";
                when x"809" => data <= "10100";
                when x"80A" => data <= "10100";
                when x"80B" => data <= "01011";
                when x"80C" => data <= "00000";
                when x"80D" => data <= "00110";
                when x"80E" => data <= "00000";
                when x"80F" => data <= "00110";
                when x"810" => data <= "00000";
                when x"811" => data <= "00110";
                when x"812" => data <= "00000";
                when x"813" => data <= "00110";
                when x"814" => data <= "00110";
                when x"815" => data <= "11100";
                when x"816" => data <= "00110";
                when x"817" => data <= "00000";
                when x"818" => data <= "10010";
                when x"819" => data <= "00000";
                when x"81A" => data <= "00110";
                when x"81B" => data <= "00000";
                when x"81C" => data <= "00000";
                when x"81D" => data <= "00000";
                when x"81E" => data <= "00110";
                when x"81F" => data <= "00000";
                when x"820" => data <= "00000";
                when x"821" => data <= "00000";
                when x"822" => data <= "00000";
                when x"823" => data <= "00110";
                when x"824" => data <= "00110";
                when x"825" => data <= "00000";
                when x"826" => data <= "00000";
                when x"827" => data <= "00000";
                when x"828" => data <= "00000";
                when x"829" => data <= "00000";
                when x"82A" => data <= "00110";
                when x"82B" => data <= "00000";
                when x"82C" => data <= "00110";
                when x"82D" => data <= "00000";
                when x"82E" => data <= "00110";
                when x"82F" => data <= "00110";
                when x"830" => data <= "01101";
                when x"831" => data <= "01101";
                when x"832" => data <= "00000";
                when x"833" => data <= "00000";
                when x"834" => data <= "00000";
                when x"835" => data <= "00000";
                when x"836" => data <= "00000";
                when x"837" => data <= "10110";
                when x"838" => data <= "00110";
                when x"839" => data <= "00000";
                when x"83A" => data <= "00000";
                when x"83B" => data <= "11010";
                when x"83C" => data <= "00000";
                when x"83D" => data <= "00110";
                when x"83E" => data <= "00110";
                when x"83F" => data <= "11001";
                when x"840" => data <= "00110";
                when x"841" => data <= "00110";
                when x"842" => data <= "10101";
                when x"843" => data <= "11111";
                when x"844" => data <= "00110";
                when x"845" => data <= "00110";
                when x"846" => data <= "00000";
                when x"847" => data <= "01111";
                when x"848" => data <= "00110";
                when x"849" => data <= "00000";
                when x"84A" => data <= "00110";
                when x"84B" => data <= "00000";
                when x"84C" => data <= "01011";
                when x"84D" => data <= "00011";
                when x"84E" => data <= "00110";
                when x"84F" => data <= "00110";
                when x"850" => data <= "10011";
                when x"851" => data <= "00000";
                when x"852" => data <= "00110";
                when x"853" => data <= "00000";
                when x"854" => data <= "00110";
                when x"855" => data <= "00000";
                when x"856" => data <= "00000";
                when x"857" => data <= "00000";
                when x"858" => data <= "00000";
                when x"859" => data <= "00110";
                when x"85A" => data <= "00010";
                when x"85B" => data <= "00000";
                when x"85C" => data <= "00000";
                when x"85D" => data <= "00000";
                when x"85E" => data <= "00001";
                when x"85F" => data <= "00000";
                when x"860" => data <= "00110";
                when x"861" => data <= "00111";
                when x"862" => data <= "00000";
                when x"863" => data <= "00110";
                when x"864" => data <= "00000";
                when x"865" => data <= "10100";
                when x"866" => data <= "00000";
                when x"867" => data <= "00110";
                when x"868" => data <= "00000";
                when x"869" => data <= "00000";
                when x"86A" => data <= "00000";
                when x"86B" => data <= "00110";
                when x"86C" => data <= "00110";
                when x"86D" => data <= "00110";
                when x"86E" => data <= "00000";
                when x"86F" => data <= "00110";
                when x"870" => data <= "00110";
                when x"871" => data <= "00110";
                when x"872" => data <= "00110";
                when x"873" => data <= "00000";
                when x"874" => data <= "01011";
                when x"875" => data <= "00000";
                when x"876" => data <= "00110";
                when x"877" => data <= "10111";
                when x"878" => data <= "00110";
                when x"879" => data <= "00110";
                when x"87A" => data <= "00000";
                when x"87B" => data <= "00110";
                when x"87C" => data <= "01101";
                when x"87D" => data <= "00000";
                when x"87E" => data <= "00000";
                when x"87F" => data <= "00000";
                when x"880" => data <= "01011";
                when x"881" => data <= "00000";
                when x"882" => data <= "10110";
                when x"883" => data <= "01100";
                when x"884" => data <= "00000";
                when x"885" => data <= "00110";
                when x"886" => data <= "00110";
                when x"887" => data <= "00000";
                when x"888" => data <= "00000";
                when x"889" => data <= "00000";
                when x"88A" => data <= "00000";
                when x"88B" => data <= "00000";
                when x"88C" => data <= "00110";
                when x"88D" => data <= "00000";
                when x"88E" => data <= "00110";
                when x"88F" => data <= "00000";
                when x"890" => data <= "00110";
                when x"891" => data <= "01101";
                when x"892" => data <= "11011";
                when x"893" => data <= "00000";
                when x"894" => data <= "00110";
                when x"895" => data <= "11101";
                when x"896" => data <= "00110";
                when x"897" => data <= "00110";
                when x"898" => data <= "00000";
                when x"899" => data <= "00110";
                when x"89A" => data <= "00110";
                when x"89B" => data <= "00110";
                when x"89C" => data <= "11000";
                when x"89D" => data <= "00110";
                when x"89E" => data <= "00110";
                when x"89F" => data <= "00110";
                when x"8A0" => data <= "00110";
                when x"8A1" => data <= "00110";
                when x"8A2" => data <= "00110";
                when x"8A3" => data <= "11001";
                when x"8A4" => data <= "00011";
                when x"8A5" => data <= "00000";
                when x"8A6" => data <= "00100";
                when x"8A7" => data <= "00110";
                when x"8A8" => data <= "00110";
                when x"8A9" => data <= "00000";
                when x"8AA" => data <= "00000";
                when x"8AB" => data <= "00110";
                when x"8AC" => data <= "00110";
                when x"8AD" => data <= "00000";
                when x"8AE" => data <= "00110";
                when x"8AF" => data <= "01011";
                when x"8B0" => data <= "00000";
                when x"8B1" => data <= "10011";
                when x"8B2" => data <= "10010";
                when x"8B3" => data <= "11110";
                when x"8B4" => data <= "00000";
                when x"8B5" => data <= "00110";
                when x"8B6" => data <= "01100";
                when x"8B7" => data <= "00000";
                when x"8B8" => data <= "11010";
                when x"8B9" => data <= "00110";
                when x"8BA" => data <= "00000";
                when x"8BB" => data <= "00000";
                when x"8BC" => data <= "00000";
                when x"8BD" => data <= "00000";
                when x"8BE" => data <= "00000";
                when x"8BF" => data <= "00110";
                when x"8C0" => data <= "00110";
                when x"8C1" => data <= "00000";
                when x"8C2" => data <= "00000";
                when x"8C3" => data <= "00000";
                when x"8C4" => data <= "00000";
                when x"8C5" => data <= "10111";
                when x"8C6" => data <= "00110";
                when x"8C7" => data <= "00000";
                when x"8C8" => data <= "00000";
                when x"8C9" => data <= "00110";
                when x"8CA" => data <= "00110";
                when x"8CB" => data <= "00110";
                when x"8CC" => data <= "00000";
                when x"8CD" => data <= "01011";
                when x"8CE" => data <= "11000";
                when x"8CF" => data <= "00000";
                when x"8D0" => data <= "00111";
                when x"8D1" => data <= "00110";
                when x"8D2" => data <= "00110";
                when x"8D3" => data <= "01000";
                when x"8D4" => data <= "00110";
                when x"8D5" => data <= "00110";
                when x"8D6" => data <= "00111";
                when x"8D7" => data <= "00110";
                when x"8D8" => data <= "00000";
                when x"8D9" => data <= "00000";
                when x"8DA" => data <= "00000";
                when x"8DB" => data <= "00000";
                when x"8DC" => data <= "00000";
                when x"8DD" => data <= "00110";
                when x"8DE" => data <= "00000";
                when x"8DF" => data <= "00110";
                when x"8E0" => data <= "00000";
                when x"8E1" => data <= "00000";
                when x"8E2" => data <= "00001";
                when x"8E3" => data <= "00000";
                when x"8E4" => data <= "00110";
                when x"8E5" => data <= "00000";
                when x"8E6" => data <= "00010";
                when x"8E7" => data <= "00000";
                when x"8E8" => data <= "00011";
                when x"8E9" => data <= "00000";
                when x"8EA" => data <= "00110";
                when x"8EB" => data <= "00000";
                when x"8EC" => data <= "00111";
                when x"8ED" => data <= "00000";
                when x"8EE" => data <= "00110";
                when x"8EF" => data <= "00000";
                when x"8F0" => data <= "00110";
                when x"8F1" => data <= "00000";
                when x"8F2" => data <= "00000";
                when x"8F3" => data <= "00000";
                when x"8F4" => data <= "00110";
                when x"8F5" => data <= "01001";
                when x"8F6" => data <= "00000";
                when x"8F7" => data <= "00110";
                when x"8F8" => data <= "00000";
                when x"8F9" => data <= "01001";
                when x"8FA" => data <= "00110";
                when x"8FB" => data <= "00000";
                when x"8FC" => data <= "00110";
                when x"8FD" => data <= "00110";
                when x"8FE" => data <= "00110";
                when x"8FF" => data <= "00110";
                when x"900" => data <= "01101";
                when x"901" => data <= "00000";
                when x"902" => data <= "00000";
                when x"903" => data <= "10110";
                when x"904" => data <= "10011";
                when x"905" => data <= "01000";
                when x"906" => data <= "00110";
                when x"907" => data <= "00110";
                when x"908" => data <= "00000";
                when x"909" => data <= "00000";
                when x"90A" => data <= "00000";
                when x"90B" => data <= "00000";
                when x"90C" => data <= "00110";
                when x"90D" => data <= "00110";
                when x"90E" => data <= "00000";
                when x"90F" => data <= "00110";
                when x"910" => data <= "01011";
                when x"911" => data <= "00110";
                when x"912" => data <= "00000";
                when x"913" => data <= "00000";
                when x"914" => data <= "00000";
                when x"915" => data <= "00110";
                when x"916" => data <= "00000";
                when x"917" => data <= "00110";
                when x"918" => data <= "00000";
                when x"919" => data <= "00000";
                when x"91A" => data <= "00110";
                when x"91B" => data <= "00100";
                when x"91C" => data <= "00000";
                when x"91D" => data <= "00000";
                when x"91E" => data <= "10011";
                when x"91F" => data <= "00110";
                when x"920" => data <= "11000";
                when x"921" => data <= "10011";
                when x"922" => data <= "00000";
                when x"923" => data <= "11101";
                when x"924" => data <= "00110";
                when x"925" => data <= "00000";
                when x"926" => data <= "00110";
                when x"927" => data <= "00110";
                when x"928" => data <= "00000";
                when x"929" => data <= "11010";
                when x"92A" => data <= "11001";
                when x"92B" => data <= "01011";
                when x"92C" => data <= "10000";
                when x"92D" => data <= "00110";
                when x"92E" => data <= "00110";
                when x"92F" => data <= "00000";
                when x"930" => data <= "00111";
                when x"931" => data <= "00000";
                when x"932" => data <= "00110";
                when x"933" => data <= "00000";
                when x"934" => data <= "00110";
                when x"935" => data <= "00110";
                when x"936" => data <= "00000";
                when x"937" => data <= "00000";
                when x"938" => data <= "00110";
                when x"939" => data <= "00101";
                when x"93A" => data <= "00000";
                when x"93B" => data <= "00110";
                when x"93C" => data <= "00110";
                when x"93D" => data <= "00000";
                when x"93E" => data <= "00000";
                when x"93F" => data <= "00110";
                when x"940" => data <= "00011";
                when x"941" => data <= "00110";
                when x"942" => data <= "10100";
                when x"943" => data <= "00000";
                when x"944" => data <= "00000";
                when x"945" => data <= "01100";
                when x"946" => data <= "00110";
                when x"947" => data <= "00100";
                when x"948" => data <= "01011";
                when x"949" => data <= "01011";
                when x"94A" => data <= "01101";
                when x"94B" => data <= "00000";
                when x"94C" => data <= "00110";
                when x"94D" => data <= "01101";
                when x"94E" => data <= "00110";
                when x"94F" => data <= "00110";
                when x"950" => data <= "00110";
                when x"951" => data <= "00000";
                when x"952" => data <= "00000";
                when x"953" => data <= "00110";
                when x"954" => data <= "00110";
                when x"955" => data <= "00000";
                when x"956" => data <= "00000";
                when x"957" => data <= "00000";
                when x"958" => data <= "00110";
                when x"959" => data <= "00110";
                when x"95A" => data <= "00000";
                when x"95B" => data <= "00000";
                when x"95C" => data <= "00000";
                when x"95D" => data <= "00000";
                when x"95E" => data <= "00110";
                when x"95F" => data <= "00000";
                when x"960" => data <= "00110";
                when x"961" => data <= "00110";
                when x"962" => data <= "00110";
                when x"963" => data <= "00110";
                when x"964" => data <= "00000";
                when x"965" => data <= "00110";
                when x"966" => data <= "00000";
                when x"967" => data <= "00000";
                when x"968" => data <= "00111";
                when x"969" => data <= "00000";
                when x"96A" => data <= "00000";
                when x"96B" => data <= "00000";
                when x"96C" => data <= "00110";
                when x"96D" => data <= "00110";
                when x"96E" => data <= "00000";
                when x"96F" => data <= "00110";
                when x"970" => data <= "10101";
                when x"971" => data <= "01011";
                when x"972" => data <= "00000";
                when x"973" => data <= "00110";
                when x"974" => data <= "00110";
                when x"975" => data <= "00000";
                when x"976" => data <= "00110";
                when x"977" => data <= "11000";
                when x"978" => data <= "00110";
                when x"979" => data <= "01010";
                when x"97A" => data <= "00110";
                when x"97B" => data <= "00000";
                when x"97C" => data <= "01101";
                when x"97D" => data <= "00000";
                when x"97E" => data <= "00000";
                when x"97F" => data <= "00110";
                when x"980" => data <= "00110";
                when x"981" => data <= "00000";
                when x"982" => data <= "00000";
                when x"983" => data <= "11001";
                when x"984" => data <= "00110";
                when x"985" => data <= "00000";
                when x"986" => data <= "00000";
                when x"987" => data <= "00110";
                when x"988" => data <= "00000";
                when x"989" => data <= "00000";
                when x"98A" => data <= "01011";
                when x"98B" => data <= "00110";
                when x"98C" => data <= "00000";
                when x"98D" => data <= "10101";
                when x"98E" => data <= "00110";
                when x"98F" => data <= "00110";
                when x"990" => data <= "00000";
                when x"991" => data <= "00000";
                when x"992" => data <= "11110";
                when x"993" => data <= "00110";
                when x"994" => data <= "00111";
                when x"995" => data <= "00110";
                when x"996" => data <= "00000";
                when x"997" => data <= "00000";
                when x"998" => data <= "00110";
                when x"999" => data <= "00000";
                when x"99A" => data <= "00000";
                when x"99B" => data <= "00000";
                when x"99C" => data <= "00000";
                when x"99D" => data <= "00110";
                when x"99E" => data <= "00110";
                when x"99F" => data <= "00000";
                when x"9A0" => data <= "00110";
                when x"9A1" => data <= "00110";
                when x"9A2" => data <= "00110";
                when x"9A3" => data <= "00000";
                when x"9A4" => data <= "00000";
                when x"9A5" => data <= "11001";
                when x"9A6" => data <= "00110";
                when x"9A7" => data <= "11011";
                when x"9A8" => data <= "00110";
                when x"9A9" => data <= "00000";
                when x"9AA" => data <= "00110";
                when x"9AB" => data <= "00110";
                when x"9AC" => data <= "11000";
                when x"9AD" => data <= "00110";
                when x"9AE" => data <= "00111";
                when x"9AF" => data <= "00110";
                when x"9B0" => data <= "11110";
                when x"9B1" => data <= "00110";
                when x"9B2" => data <= "00110";
                when x"9B3" => data <= "00111";
                when x"9B4" => data <= "00110";
                when x"9B5" => data <= "01110";
                when x"9B6" => data <= "01101";
                when x"9B7" => data <= "00110";
                when x"9B8" => data <= "00110";
                when x"9B9" => data <= "01101";
                when x"9BA" => data <= "00000";
                when x"9BB" => data <= "11100";
                when x"9BC" => data <= "00110";
                when x"9BD" => data <= "00110";
                when x"9BE" => data <= "00110";
                when x"9BF" => data <= "00110";
                when x"9C0" => data <= "00000";
                when x"9C1" => data <= "00000";
                when x"9C2" => data <= "00110";
                when x"9C3" => data <= "00011";
                when x"9C4" => data <= "01101";
                when x"9C5" => data <= "01010";
                when x"9C6" => data <= "00000";
                when x"9C7" => data <= "00000";
                when x"9C8" => data <= "00000";
                when x"9C9" => data <= "00110";
                when x"9CA" => data <= "00110";
                when x"9CB" => data <= "00000";
                when x"9CC" => data <= "00000";
                when x"9CD" => data <= "00110";
                when x"9CE" => data <= "00110";
                when x"9CF" => data <= "00110";
                when x"9D0" => data <= "00110";
                when x"9D1" => data <= "01110";
                when x"9D2" => data <= "00000";
                when x"9D3" => data <= "00000";
                when x"9D4" => data <= "00000";
                when x"9D5" => data <= "00110";
                when x"9D6" => data <= "00000";
                when x"9D7" => data <= "00110";
                when x"9D8" => data <= "00000";
                when x"9D9" => data <= "00000";
                when x"9DA" => data <= "00000";
                when x"9DB" => data <= "00000";
                when x"9DC" => data <= "00000";
                when x"9DD" => data <= "00110";
                when x"9DE" => data <= "00110";
                when x"9DF" => data <= "00110";
                when x"9E0" => data <= "01011";
                when x"9E1" => data <= "00000";
                when x"9E2" => data <= "01001";
                when x"9E3" => data <= "00110";
                when x"9E4" => data <= "00000";
                when x"9E5" => data <= "00000";
                when x"9E6" => data <= "00000";
                when x"9E7" => data <= "00110";
                when x"9E8" => data <= "00000";
                when x"9E9" => data <= "00000";
                when x"9EA" => data <= "00000";
                when x"9EB" => data <= "00110";
                when x"9EC" => data <= "00110";
                when x"9ED" => data <= "00000";
                when x"9EE" => data <= "00000";
                when x"9EF" => data <= "00110";
                when x"9F0" => data <= "00000";
                when x"9F1" => data <= "01101";
                when x"9F2" => data <= "00000";
                when x"9F3" => data <= "00000";
                when x"9F4" => data <= "00000";
                when x"9F5" => data <= "00000";
                when x"9F6" => data <= "00000";
                when x"9F7" => data <= "00110";
                when x"9F8" => data <= "00110";
                when x"9F9" => data <= "00000";
                when x"9FA" => data <= "11001";
                when x"9FB" => data <= "00000";
                when x"9FC" => data <= "00110";
                when x"9FD" => data <= "11001";
                when x"9FE" => data <= "00110";
                when x"9FF" => data <= "00000";
                when x"A00" => data <= "00110";
                when x"A01" => data <= "00000";
                when x"A02" => data <= "00000";
                when x"A03" => data <= "00110";
                when x"A04" => data <= "00110";
                when x"A05" => data <= "00111";
                when x"A06" => data <= "00110";
                when x"A07" => data <= "01101";
                when x"A08" => data <= "00110";
                when x"A09" => data <= "00110";
                when x"A0A" => data <= "00000";
                when x"A0B" => data <= "00110";
                when x"A0C" => data <= "00110";
                when x"A0D" => data <= "00000";
                when x"A0E" => data <= "00000";
                when x"A0F" => data <= "00000";
                when x"A10" => data <= "00000";
                when x"A11" => data <= "00110";
                when x"A12" => data <= "00110";
                when x"A13" => data <= "10100";
                when x"A14" => data <= "00000";
                when x"A15" => data <= "00000";
                when x"A16" => data <= "00000";
                when x"A17" => data <= "00000";
                when x"A18" => data <= "10111";
                when x"A19" => data <= "00000";
                when x"A1A" => data <= "01011";
                when x"A1B" => data <= "00010";
                when x"A1C" => data <= "00101";
                when x"A1D" => data <= "00000";
                when x"A1E" => data <= "00110";
                when x"A1F" => data <= "00110";
                when x"A20" => data <= "11100";
                when x"A21" => data <= "00101";
                when x"A22" => data <= "11111";
                when x"A23" => data <= "00000";
                when x"A24" => data <= "00000";
                when x"A25" => data <= "00110";
                when x"A26" => data <= "10100";
                when x"A27" => data <= "00110";
                when x"A28" => data <= "00110";
                when x"A29" => data <= "00000";
                when x"A2A" => data <= "00110";
                when x"A2B" => data <= "00110";
                when x"A2C" => data <= "00110";
                when x"A2D" => data <= "00110";
                when x"A2E" => data <= "00110";
                when x"A2F" => data <= "00000";
                when x"A30" => data <= "00000";
                when x"A31" => data <= "00110";
                when x"A32" => data <= "01011";
                when x"A33" => data <= "00000";
                when x"A34" => data <= "00000";
                when x"A35" => data <= "00110";
                when x"A36" => data <= "00000";
                when x"A37" => data <= "00000";
                when x"A38" => data <= "00110";
                when x"A39" => data <= "00000";
                when x"A3A" => data <= "01011";
                when x"A3B" => data <= "11001";
                when x"A3C" => data <= "00110";
                when x"A3D" => data <= "00000";
                when x"A3E" => data <= "00000";
                when x"A3F" => data <= "11001";
                when x"A40" => data <= "00000";
                when x"A41" => data <= "00000";
                when x"A42" => data <= "00000";
                when x"A43" => data <= "00110";
                when x"A44" => data <= "10110";
                when x"A45" => data <= "00000";
                when x"A46" => data <= "00110";
                when x"A47" => data <= "00110";
                when x"A48" => data <= "00000";
                when x"A49" => data <= "10111";
                when x"A4A" => data <= "00000";
                when x"A4B" => data <= "00000";
                when x"A4C" => data <= "00110";
                when x"A4D" => data <= "00110";
                when x"A4E" => data <= "00000";
                when x"A4F" => data <= "00110";
                when x"A50" => data <= "00000";
                when x"A51" => data <= "00110";
                when x"A52" => data <= "00000";
                when x"A53" => data <= "00000";
                when x"A54" => data <= "10011";
                when x"A55" => data <= "10011";
                when x"A56" => data <= "00000";
                when x"A57" => data <= "00000";
                when x"A58" => data <= "00110";
                when x"A59" => data <= "00110";
                when x"A5A" => data <= "00110";
                when x"A5B" => data <= "00000";
                when x"A5C" => data <= "01101";
                when x"A5D" => data <= "00000";
                when x"A5E" => data <= "00000";
                when x"A5F" => data <= "00000";
                when x"A60" => data <= "01101";
                when x"A61" => data <= "00101";
                when x"A62" => data <= "00110";
                when x"A63" => data <= "00110";
                when x"A64" => data <= "00000";
                when x"A65" => data <= "00000";
                when x"A66" => data <= "01011";
                when x"A67" => data <= "00000";
                when x"A68" => data <= "11010";
                when x"A69" => data <= "00110";
                when x"A6A" => data <= "00001";
                when x"A6B" => data <= "11010";
                when x"A6C" => data <= "01100";
                when x"A6D" => data <= "01100";
                when x"A6E" => data <= "00000";
                when x"A6F" => data <= "00010";
                when x"A70" => data <= "00000";
                when x"A71" => data <= "11111";
                when x"A72" => data <= "00000";
                when x"A73" => data <= "00110";
                when x"A74" => data <= "00000";
                when x"A75" => data <= "00000";
                when x"A76" => data <= "00000";
                when x"A77" => data <= "00000";
                when x"A78" => data <= "00110";
                when x"A79" => data <= "00110";
                when x"A7A" => data <= "00000";
                when x"A7B" => data <= "00000";
                when x"A7C" => data <= "00000";
                when x"A7D" => data <= "00110";
                when x"A7E" => data <= "00000";
                when x"A7F" => data <= "00110";
                when x"A80" => data <= "00110";
                when x"A81" => data <= "01101";
                when x"A82" => data <= "01010";
                when x"A83" => data <= "00000";
                when x"A84" => data <= "11000";
                when x"A85" => data <= "01101";
                when x"A86" => data <= "00110";
                when x"A87" => data <= "00110";
                when x"A88" => data <= "00000";
                when x"A89" => data <= "10111";
                when x"A8A" => data <= "00000";
                when x"A8B" => data <= "00000";
                when x"A8C" => data <= "11001";
                when x"A8D" => data <= "10010";
                when x"A8E" => data <= "01101";
                when x"A8F" => data <= "00000";
                when x"A90" => data <= "00110";
                when x"A91" => data <= "00000";
                when x"A92" => data <= "00110";
                when x"A93" => data <= "01000";
                when x"A94" => data <= "00110";
                when x"A95" => data <= "00110";
                when x"A96" => data <= "11100";
                when x"A97" => data <= "00011";
                when x"A98" => data <= "11110";
                when x"A99" => data <= "00000";
                when x"A9A" => data <= "00000";
                when x"A9B" => data <= "00000";
                when x"A9C" => data <= "00000";
                when x"A9D" => data <= "00000";
                when x"A9E" => data <= "00110";
                when x"A9F" => data <= "00110";
                when x"AA0" => data <= "00110";
                when x"AA1" => data <= "00000";
                when x"AA2" => data <= "01110";
                when x"AA3" => data <= "11001";
                when x"AA4" => data <= "00000";
                when x"AA5" => data <= "10110";
                when x"AA6" => data <= "00000";
                when x"AA7" => data <= "00110";
                when x"AA8" => data <= "00110";
                when x"AA9" => data <= "00110";
                when x"AAA" => data <= "11110";
                when x"AAB" => data <= "00000";
                when x"AAC" => data <= "00111";
                when x"AAD" => data <= "01001";
                when x"AAE" => data <= "00110";
                when x"AAF" => data <= "00110";
                when x"AB0" => data <= "00110";
                when x"AB1" => data <= "00110";
                when x"AB2" => data <= "01100";
                when x"AB3" => data <= "11100";
                when x"AB4" => data <= "00110";
                when x"AB5" => data <= "10100";
                when x"AB6" => data <= "01110";
                when x"AB7" => data <= "00000";
                when x"AB8" => data <= "00110";
                when x"AB9" => data <= "00110";
                when x"ABA" => data <= "00000";
                when x"ABB" => data <= "00110";
                when x"ABC" => data <= "00000";
                when x"ABD" => data <= "01101";
                when x"ABE" => data <= "00000";
                when x"ABF" => data <= "00000";
                when x"AC0" => data <= "00100";
                when x"AC1" => data <= "00000";
                when x"AC2" => data <= "00110";
                when x"AC3" => data <= "00000";
                when x"AC4" => data <= "00110";
                when x"AC5" => data <= "00110";
                when x"AC6" => data <= "00110";
                when x"AC7" => data <= "01010";
                when x"AC8" => data <= "00000";
                when x"AC9" => data <= "00000";
                when x"ACA" => data <= "00000";
                when x"ACB" => data <= "00110";
                when x"ACC" => data <= "01000";
                when x"ACD" => data <= "00000";
                when x"ACE" => data <= "00110";
                when x"ACF" => data <= "01101";
                when x"AD0" => data <= "00110";
                when x"AD1" => data <= "00110";
                when x"AD2" => data <= "00000";
                when x"AD3" => data <= "00000";
                when x"AD4" => data <= "00110";
                when x"AD5" => data <= "10011";
                when x"AD6" => data <= "00000";
                when x"AD7" => data <= "00110";
                when x"AD8" => data <= "00000";
                when x"AD9" => data <= "00110";
                when x"ADA" => data <= "00000";
                when x"ADB" => data <= "00000";
                when x"ADC" => data <= "00000";
                when x"ADD" => data <= "00110";
                when x"ADE" => data <= "00000";
                when x"ADF" => data <= "10000";
                when x"AE0" => data <= "00000";
                when x"AE1" => data <= "01010";
                when x"AE2" => data <= "00000";
                when x"AE3" => data <= "00000";
                when x"AE4" => data <= "00110";
                when x"AE5" => data <= "11000";
                when x"AE6" => data <= "00110";
                when x"AE7" => data <= "10011";
                when x"AE8" => data <= "11111";
                when x"AE9" => data <= "00110";
                when x"AEA" => data <= "00110";
                when x"AEB" => data <= "00110";
                when x"AEC" => data <= "00000";
                when x"AED" => data <= "00110";
                when x"AEE" => data <= "00110";
                when x"AEF" => data <= "00110";
                when x"AF0" => data <= "00110";
                when x"AF1" => data <= "10101";
                when x"AF2" => data <= "00110";
                when x"AF3" => data <= "00000";
                when x"AF4" => data <= "00000";
                when x"AF5" => data <= "00000";
                when x"AF6" => data <= "00110";
                when x"AF7" => data <= "00110";
                when x"AF8" => data <= "00000";
                when x"AF9" => data <= "00000";
                when x"AFA" => data <= "00011";
                when x"AFB" => data <= "00000";
                when x"AFC" => data <= "00000";
                when x"AFD" => data <= "00110";
                when x"AFE" => data <= "00000";
                when x"AFF" => data <= "00110";
                when x"B00" => data <= "00000";
                when x"B01" => data <= "00110";
                when x"B02" => data <= "00110";
                when x"B03" => data <= "00110";
                when x"B04" => data <= "00110";
                when x"B05" => data <= "11101";
                when x"B06" => data <= "00000";
                when x"B07" => data <= "10011";
                when x"B08" => data <= "00000";
                when x"B09" => data <= "00110";
                when x"B0A" => data <= "01001";
                when x"B0B" => data <= "00110";
                when x"B0C" => data <= "00110";
                when x"B0D" => data <= "00000";
                when x"B0E" => data <= "00001";
                when x"B0F" => data <= "00000";
                when x"B10" => data <= "00000";
                when x"B11" => data <= "11001";
                when x"B12" => data <= "00110";
                when x"B13" => data <= "00110";
                when x"B14" => data <= "00110";
                when x"B15" => data <= "00000";
                when x"B16" => data <= "00110";
                when x"B17" => data <= "10010";
                when x"B18" => data <= "00110";
                when x"B19" => data <= "00000";
                when x"B1A" => data <= "00111";
                when x"B1B" => data <= "00000";
                when x"B1C" => data <= "00000";
                when x"B1D" => data <= "00110";
                when x"B1E" => data <= "00110";
                when x"B1F" => data <= "00110";
                when x"B20" => data <= "00000";
                when x"B21" => data <= "10000";
                when x"B22" => data <= "00000";
                when x"B23" => data <= "00110";
                when x"B24" => data <= "00000";
                when x"B25" => data <= "00000";
                when x"B26" => data <= "11001";
                when x"B27" => data <= "00000";
                when x"B28" => data <= "00000";
                when x"B29" => data <= "10100";
                when x"B2A" => data <= "00110";
                when x"B2B" => data <= "00110";
                when x"B2C" => data <= "00000";
                when x"B2D" => data <= "00110";
                when x"B2E" => data <= "00000";
                when x"B2F" => data <= "00000";
                when x"B30" => data <= "11110";
                when x"B31" => data <= "00000";
                when x"B32" => data <= "00110";
                when x"B33" => data <= "00000";
                when x"B34" => data <= "00110";
                when x"B35" => data <= "00110";
                when x"B36" => data <= "00110";
                when x"B37" => data <= "00110";
                when x"B38" => data <= "00110";
                when x"B39" => data <= "00000";
                when x"B3A" => data <= "00000";
                when x"B3B" => data <= "00000";
                when x"B3C" => data <= "00000";
                when x"B3D" => data <= "00110";
                when x"B3E" => data <= "00000";
                when x"B3F" => data <= "00000";
                when x"B40" => data <= "00101";
                when x"B41" => data <= "00000";
                when x"B42" => data <= "00110";
                when x"B43" => data <= "00110";
                when x"B44" => data <= "00000";
                when x"B45" => data <= "00000";
                when x"B46" => data <= "00110";
                when x"B47" => data <= "00000";
                when x"B48" => data <= "10110";
                when x"B49" => data <= "00000";
                when x"B4A" => data <= "00000";
                when x"B4B" => data <= "00110";
                when x"B4C" => data <= "00000";
                when x"B4D" => data <= "00110";
                when x"B4E" => data <= "01101";
                when x"B4F" => data <= "00000";
                when x"B50" => data <= "10010";
                when x"B51" => data <= "00000";
                when x"B52" => data <= "00110";
                when x"B53" => data <= "00000";
                when x"B54" => data <= "00101";
                when x"B55" => data <= "00111";
                when x"B56" => data <= "00110";
                when x"B57" => data <= "00110";
                when x"B58" => data <= "00110";
                when x"B59" => data <= "00110";
                when x"B5A" => data <= "00110";
                when x"B5B" => data <= "00000";
                when x"B5C" => data <= "00000";
                when x"B5D" => data <= "00110";
                when x"B5E" => data <= "00000";
                when x"B5F" => data <= "00110";
                when x"B60" => data <= "00000";
                when x"B61" => data <= "00000";
                when x"B62" => data <= "00110";
                when x"B63" => data <= "10111";
                when x"B64" => data <= "00000";
                when x"B65" => data <= "00000";
                when x"B66" => data <= "01101";
                when x"B67" => data <= "00000";
                when x"B68" => data <= "00110";
                when x"B69" => data <= "00000";
                when x"B6A" => data <= "00110";
                when x"B6B" => data <= "00000";
                when x"B6C" => data <= "00000";
                when x"B6D" => data <= "00001";
                when x"B6E" => data <= "00000";
                when x"B6F" => data <= "00000";
                when x"B70" => data <= "00110";
                when x"B71" => data <= "01101";
                when x"B72" => data <= "00000";
                when x"B73" => data <= "00000";
                when x"B74" => data <= "00000";
                when x"B75" => data <= "00000";
                when x"B76" => data <= "11111";
                when x"B77" => data <= "00110";
                when x"B78" => data <= "00000";
                when x"B79" => data <= "00000";
                when x"B7A" => data <= "00110";
                when x"B7B" => data <= "00010";
                when x"B7C" => data <= "11011";
                when x"B7D" => data <= "00000";
                when x"B7E" => data <= "00110";
                when x"B7F" => data <= "00110";
                when x"B80" => data <= "01011";
                when x"B81" => data <= "00000";
                when x"B82" => data <= "00110";
                when x"B83" => data <= "00000";
                when x"B84" => data <= "00000";
                when x"B85" => data <= "11001";
                when x"B86" => data <= "00000";
                when x"B87" => data <= "00110";
                when x"B88" => data <= "00110";
                when x"B89" => data <= "01000";
                when x"B8A" => data <= "00000";
                when x"B8B" => data <= "00110";
                when x"B8C" => data <= "00000";
                when x"B8D" => data <= "01011";
                when x"B8E" => data <= "00110";
                when x"B8F" => data <= "00000";
                when x"B90" => data <= "00000";
                when x"B91" => data <= "01000";
                when x"B92" => data <= "01110";
                when x"B93" => data <= "10010";
                when x"B94" => data <= "00000";
                when x"B95" => data <= "00001";
                when x"B96" => data <= "00110";
                when x"B97" => data <= "00000";
                when x"B98" => data <= "10111";
                when x"B99" => data <= "00110";
                when x"B9A" => data <= "00000";
                when x"B9B" => data <= "00110";
                when x"B9C" => data <= "00000";
                when x"B9D" => data <= "00000";
                when x"B9E" => data <= "00000";
                when x"B9F" => data <= "00000";
                when x"BA0" => data <= "00000";
                when x"BA1" => data <= "01101";
                when x"BA2" => data <= "00110";
                when x"BA3" => data <= "00110";
                when x"BA4" => data <= "00110";
                when x"BA5" => data <= "00000";
                when x"BA6" => data <= "00110";
                when x"BA7" => data <= "00000";
                when x"BA8" => data <= "00110";
                when x"BA9" => data <= "01010";
                when x"BAA" => data <= "00110";
                when x"BAB" => data <= "00011";
                when x"BAC" => data <= "00000";
                when x"BAD" => data <= "00000";
                when x"BAE" => data <= "01100";
                when x"BAF" => data <= "00000";
                when x"BB0" => data <= "00110";
                when x"BB1" => data <= "00000";
                when x"BB2" => data <= "01010";
                when x"BB3" => data <= "00000";
                when x"BB4" => data <= "00110";
                when x"BB5" => data <= "00000";
                when x"BB6" => data <= "00000";
                when x"BB7" => data <= "01001";
                when x"BB8" => data <= "00110";
                when x"BB9" => data <= "00110";
                when x"BBA" => data <= "00110";
                when x"BBB" => data <= "00000";
                when x"BBC" => data <= "10111";
                when x"BBD" => data <= "10000";
                when x"BBE" => data <= "00000";
                when x"BBF" => data <= "00000";
                when x"BC0" => data <= "00110";
                when x"BC1" => data <= "00110";
                when x"BC2" => data <= "00110";
                when x"BC3" => data <= "00000";
                when x"BC4" => data <= "00000";
                when x"BC5" => data <= "00110";
                when x"BC6" => data <= "00110";
                when x"BC7" => data <= "00000";
                when x"BC8" => data <= "00000";
                when x"BC9" => data <= "00110";
                when x"BCA" => data <= "11111";
                when x"BCB" => data <= "00110";
                when x"BCC" => data <= "00000";
                when x"BCD" => data <= "00000";
                when x"BCE" => data <= "00000";
                when x"BCF" => data <= "00110";
                when x"BD0" => data <= "00110";
                when x"BD1" => data <= "01101";
                when x"BD2" => data <= "11111";
                when x"BD3" => data <= "00100";
                when x"BD4" => data <= "00110";
                when x"BD5" => data <= "11111";
                when x"BD6" => data <= "01001";
                when x"BD7" => data <= "00000";
                when x"BD8" => data <= "10011";
                when x"BD9" => data <= "00000";
                when x"BDA" => data <= "00000";
                when x"BDB" => data <= "11111";
                when x"BDC" => data <= "00110";
                when x"BDD" => data <= "00000";
                when x"BDE" => data <= "00111";
                when x"BDF" => data <= "01011";
                when x"BE0" => data <= "00110";
                when x"BE1" => data <= "00000";
                when x"BE2" => data <= "11111";
                when x"BE3" => data <= "00110";
                when x"BE4" => data <= "00000";
                when x"BE5" => data <= "00110";
                when x"BE6" => data <= "00000";
                when x"BE7" => data <= "00110";
                when x"BE8" => data <= "00110";
                when x"BE9" => data <= "11111";
                when x"BEA" => data <= "00000";
                when x"BEB" => data <= "00110";
                when x"BEC" => data <= "00110";
                when x"BED" => data <= "00000";
                when x"BEE" => data <= "00000";
                when x"BEF" => data <= "00000";
                when x"BF0" => data <= "00110";
                when x"BF1" => data <= "11111";
                when x"BF2" => data <= "00110";
                when x"BF3" => data <= "01111";
                when x"BF4" => data <= "00001";
                when x"BF5" => data <= "00000";
                when x"BF6" => data <= "00110";
                when x"BF7" => data <= "11111";
                when x"BF8" => data <= "11000";
                when x"BF9" => data <= "00000";
                when x"BFA" => data <= "00000";
                when x"BFB" => data <= "00110";
                when x"BFC" => data <= "00110";
                when x"BFD" => data <= "00110";
                when x"BFE" => data <= "00110";
                when x"BFF" => data <= "10001";
                when x"C00" => data <= "00000";
                when x"C01" => data <= "00000";
                when x"C02" => data <= "00110";
                when x"C03" => data <= "10100";
                when x"C04" => data <= "00110";
                when x"C05" => data <= "00000";
                when x"C06" => data <= "00110";
                when x"C07" => data <= "00110";
                when x"C08" => data <= "10001";
                when x"C09" => data <= "00000";
                when x"C0A" => data <= "00110";
                when x"C0B" => data <= "10110";
                when x"C0C" => data <= "01011";
                when x"C0D" => data <= "10000";
                when x"C0E" => data <= "00000";
                when x"C0F" => data <= "00110";
                when x"C10" => data <= "00000";
                when x"C11" => data <= "00110";
                when x"C12" => data <= "00000";
                when x"C13" => data <= "00001";
                when x"C14" => data <= "10010";
                when x"C15" => data <= "00001";
                when x"C16" => data <= "10101";
                when x"C17" => data <= "00000";
                when x"C18" => data <= "00110";
                when x"C19" => data <= "00000";
                when x"C1A" => data <= "00110";
                when x"C1B" => data <= "00110";
                when x"C1C" => data <= "00000";
                when x"C1D" => data <= "00000";
                when x"C1E" => data <= "00110";
                when x"C1F" => data <= "10111";
                when x"C20" => data <= "11010";
                when x"C21" => data <= "00110";
                when x"C22" => data <= "00100";
                when x"C23" => data <= "00000";
                when x"C24" => data <= "00000";
                when x"C25" => data <= "11111";
                when x"C26" => data <= "00110";
                when x"C27" => data <= "00110";
                when x"C28" => data <= "00110";
                when x"C29" => data <= "00110";
                when x"C2A" => data <= "00110";
                when x"C2B" => data <= "00000";
                when x"C2C" => data <= "00000";
                when x"C2D" => data <= "00110";
                when x"C2E" => data <= "00110";
                when x"C2F" => data <= "11001";
                when x"C30" => data <= "00110";
                when x"C31" => data <= "00110";
                when x"C32" => data <= "00110";
                when x"C33" => data <= "01111";
                when x"C34" => data <= "10001";
                when x"C35" => data <= "00110";
                when x"C36" => data <= "00000";
                when x"C37" => data <= "00000";
                when x"C38" => data <= "00000";
                when x"C39" => data <= "00000";
                when x"C3A" => data <= "00110";
                when x"C3B" => data <= "00110";
                when x"C3C" => data <= "00110";
                when x"C3D" => data <= "00000";
                when x"C3E" => data <= "00110";
                when x"C3F" => data <= "11100";
                when x"C40" => data <= "00000";
                when x"C41" => data <= "00110";
                when x"C42" => data <= "00000";
                when x"C43" => data <= "00000";
                when x"C44" => data <= "00000";
                when x"C45" => data <= "11001";
                when x"C46" => data <= "00110";
                when x"C47" => data <= "11000";
                when x"C48" => data <= "00110";
                when x"C49" => data <= "00000";
                when x"C4A" => data <= "01010";
                when x"C4B" => data <= "00000";
                when x"C4C" => data <= "00110";
                when x"C4D" => data <= "00000";
                when x"C4E" => data <= "00000";
                when x"C4F" => data <= "00111";
                when x"C50" => data <= "00110";
                when x"C51" => data <= "00000";
                when x"C52" => data <= "00000";
                when x"C53" => data <= "00110";
                when x"C54" => data <= "00110";
                when x"C55" => data <= "00000";
                when x"C56" => data <= "00110";
                when x"C57" => data <= "00110";
                when x"C58" => data <= "01011";
                when x"C59" => data <= "00110";
                when x"C5A" => data <= "00000";
                when x"C5B" => data <= "00110";
                when x"C5C" => data <= "00000";
                when x"C5D" => data <= "00000";
                when x"C5E" => data <= "00000";
                when x"C5F" => data <= "11111";
                when x"C60" => data <= "00110";
                when x"C61" => data <= "01101";
                when x"C62" => data <= "00000";
                when x"C63" => data <= "00110";
                when x"C64" => data <= "00000";
                when x"C65" => data <= "00110";
                when x"C66" => data <= "00000";
                when x"C67" => data <= "00000";
                when x"C68" => data <= "10011";
                when x"C69" => data <= "01011";
                when x"C6A" => data <= "00110";
                when x"C6B" => data <= "00000";
                when x"C6C" => data <= "00000";
                when x"C6D" => data <= "00000";
                when x"C6E" => data <= "00111";
                when x"C6F" => data <= "00000";
                when x"C70" => data <= "00000";
                when x"C71" => data <= "00110";
                when x"C72" => data <= "00110";
                when x"C73" => data <= "00110";
                when x"C74" => data <= "00000";
                when x"C75" => data <= "01101";
                when x"C76" => data <= "00110";
                when x"C77" => data <= "00000";
                when x"C78" => data <= "00110";
                when x"C79" => data <= "00110";
                when x"C7A" => data <= "11010";
                when x"C7B" => data <= "00110";
                when x"C7C" => data <= "11110";
                when x"C7D" => data <= "00000";
                when x"C7E" => data <= "00000";
                when x"C7F" => data <= "10010";
                when x"C80" => data <= "00110";
                when x"C81" => data <= "00110";
                when x"C82" => data <= "00000";
                when x"C83" => data <= "00000";
                when x"C84" => data <= "00000";
                when x"C85" => data <= "00000";
                when x"C86" => data <= "00000";
                when x"C87" => data <= "00110";
                when x"C88" => data <= "00000";
                when x"C89" => data <= "00000";
                when x"C8A" => data <= "00000";
                when x"C8B" => data <= "00110";
                when x"C8C" => data <= "00000";
                when x"C8D" => data <= "00000";
                when x"C8E" => data <= "00000";
                when x"C8F" => data <= "00000";
                when x"C90" => data <= "00110";
                when x"C91" => data <= "00000";
                when x"C92" => data <= "00000";
                when x"C93" => data <= "00110";
                when x"C94" => data <= "00000";
                when x"C95" => data <= "00110";
                when x"C96" => data <= "00000";
                when x"C97" => data <= "10110";
                when x"C98" => data <= "00110";
                when x"C99" => data <= "00110";
                when x"C9A" => data <= "10110";
                when x"C9B" => data <= "00000";
                when x"C9C" => data <= "00000";
                when x"C9D" => data <= "00000";
                when x"C9E" => data <= "00110";
                when x"C9F" => data <= "00110";
                when x"CA0" => data <= "00000";
                when x"CA1" => data <= "00110";
                when x"CA2" => data <= "00000";
                when x"CA3" => data <= "00000";
                when x"CA4" => data <= "01011";
                when x"CA5" => data <= "00110";
                when x"CA6" => data <= "00110";
                when x"CA7" => data <= "00110";
                when x"CA8" => data <= "00000";
                when x"CA9" => data <= "00110";
                when x"CAA" => data <= "01011";
                when x"CAB" => data <= "00110";
                when x"CAC" => data <= "00110";
                when x"CAD" => data <= "01010";
                when x"CAE" => data <= "00111";
                when x"CAF" => data <= "00000";
                when x"CB0" => data <= "00110";
                when x"CB1" => data <= "00000";
                when x"CB2" => data <= "00110";
                when x"CB3" => data <= "00000";
                when x"CB4" => data <= "10011";
                when x"CB5" => data <= "00110";
                when x"CB6" => data <= "00000";
                when x"CB7" => data <= "00000";
                when x"CB8" => data <= "00110";
                when x"CB9" => data <= "00110";
                when x"CBA" => data <= "00000";
                when x"CBB" => data <= "00000";
                when x"CBC" => data <= "00000";
                when x"CBD" => data <= "00110";
                when x"CBE" => data <= "00110";
                when x"CBF" => data <= "11101";
                when x"CC0" => data <= "00000";
                when x"CC1" => data <= "00110";
                when x"CC2" => data <= "00000";
                when x"CC3" => data <= "00000";
                when x"CC4" => data <= "01110";
                when x"CC5" => data <= "00110";
                when x"CC6" => data <= "10000";
                when x"CC7" => data <= "00000";
                when x"CC8" => data <= "00110";
                when x"CC9" => data <= "00110";
                when x"CCA" => data <= "00000";
                when x"CCB" => data <= "00000";
                when x"CCC" => data <= "00110";
                when x"CCD" => data <= "00000";
                when x"CCE" => data <= "00011";
                when x"CCF" => data <= "00000";
                when x"CD0" => data <= "00110";
                when x"CD1" => data <= "00110";
                when x"CD2" => data <= "00000";
                when x"CD3" => data <= "00110";
                when x"CD4" => data <= "00110";
                when x"CD5" => data <= "11001";
                when x"CD6" => data <= "00000";
                when x"CD7" => data <= "00000";
                when x"CD8" => data <= "00110";
                when x"CD9" => data <= "00110";
                when x"CDA" => data <= "00110";
                when x"CDB" => data <= "00110";
                when x"CDC" => data <= "00000";
                when x"CDD" => data <= "00000";
                when x"CDE" => data <= "00110";
                when x"CDF" => data <= "00000";
                when x"CE0" => data <= "11111";
                when x"CE1" => data <= "00000";
                when x"CE2" => data <= "00000";
                when x"CE3" => data <= "00110";
                when x"CE4" => data <= "00000";
                when x"CE5" => data <= "11100";
                when x"CE6" => data <= "11010";
                when x"CE7" => data <= "00000";
                when x"CE8" => data <= "00000";
                when x"CE9" => data <= "01101";
                when x"CEA" => data <= "00000";
                when x"CEB" => data <= "00000";
                when x"CEC" => data <= "00000";
                when x"CED" => data <= "00000";
                when x"CEE" => data <= "11010";
                when x"CEF" => data <= "00110";
                when x"CF0" => data <= "01101";
                when x"CF1" => data <= "00000";
                when x"CF2" => data <= "00000";
                when x"CF3" => data <= "00000";
                when x"CF4" => data <= "00000";
                when x"CF5" => data <= "00110";
                when x"CF6" => data <= "00000";
                when x"CF7" => data <= "10101";
                when x"CF8" => data <= "00110";
                when x"CF9" => data <= "00000";
                when x"CFA" => data <= "00000";
                when x"CFB" => data <= "01111";
                when x"CFC" => data <= "00000";
                when x"CFD" => data <= "11000";
                when x"CFE" => data <= "00110";
                when x"CFF" => data <= "00000";
                when x"D00" => data <= "00000";
                when x"D01" => data <= "00011";
                when x"D02" => data <= "00000";
                when x"D03" => data <= "00000";
                when x"D04" => data <= "00000";
                when x"D05" => data <= "01010";
                when x"D06" => data <= "10101";
                when x"D07" => data <= "10001";
                when x"D08" => data <= "00110";
                when x"D09" => data <= "00110";
                when x"D0A" => data <= "00000";
                when x"D0B" => data <= "00000";
                when x"D0C" => data <= "10011";
                when x"D0D" => data <= "00110";
                when x"D0E" => data <= "00000";
                when x"D0F" => data <= "10000";
                when x"D10" => data <= "00110";
                when x"D11" => data <= "00000";
                when x"D12" => data <= "00110";
                when x"D13" => data <= "01101";
                when x"D14" => data <= "00110";
                when x"D15" => data <= "00000";
                when x"D16" => data <= "00110";
                when x"D17" => data <= "00110";
                when x"D18" => data <= "00110";
                when x"D19" => data <= "10100";
                when x"D1A" => data <= "00110";
                when x"D1B" => data <= "00110";
                when x"D1C" => data <= "01010";
                when x"D1D" => data <= "00110";
                when x"D1E" => data <= "00000";
                when x"D1F" => data <= "00000";
                when x"D20" => data <= "00000";
                when x"D21" => data <= "00000";
                when x"D22" => data <= "00110";
                when x"D23" => data <= "10111";
                when x"D24" => data <= "01101";
                when x"D25" => data <= "00000";
                when x"D26" => data <= "00110";
                when x"D27" => data <= "00110";
                when x"D28" => data <= "00110";
                when x"D29" => data <= "10001";
                when x"D2A" => data <= "00110";
                when x"D2B" => data <= "00110";
                when x"D2C" => data <= "00000";
                when x"D2D" => data <= "01101";
                when x"D2E" => data <= "00100";
                when x"D2F" => data <= "00010";
                when x"D30" => data <= "00110";
                when x"D31" => data <= "00000";
                when x"D32" => data <= "00110";
                when x"D33" => data <= "01011";
                when x"D34" => data <= "00110";
                when x"D35" => data <= "00110";
                when x"D36" => data <= "00110";
                when x"D37" => data <= "00000";
                when x"D38" => data <= "00000";
                when x"D39" => data <= "00110";
                when x"D3A" => data <= "01001";
                when x"D3B" => data <= "10000";
                when x"D3C" => data <= "00110";
                when x"D3D" => data <= "10100";
                when x"D3E" => data <= "11111";
                when x"D3F" => data <= "00011";
                when x"D40" => data <= "00110";
                when x"D41" => data <= "00000";
                when x"D42" => data <= "00000";
                when x"D43" => data <= "00001";
                when x"D44" => data <= "00110";
                when x"D45" => data <= "00000";
                when x"D46" => data <= "00000";
                when x"D47" => data <= "00110";
                when x"D48" => data <= "00010";
                when x"D49" => data <= "00110";
                when x"D4A" => data <= "00000";
                when x"D4B" => data <= "00000";
                when x"D4C" => data <= "01101";
                when x"D4D" => data <= "00101";
                when x"D4E" => data <= "01110";
                when x"D4F" => data <= "00110";
                when x"D50" => data <= "00110";
                when x"D51" => data <= "00000";
                when x"D52" => data <= "00111";
                when x"D53" => data <= "00000";
                when x"D54" => data <= "00000";
                when x"D55" => data <= "00000";
                when x"D56" => data <= "00000";
                when x"D57" => data <= "01111";
                when x"D58" => data <= "10101";
                when x"D59" => data <= "00000";
                when x"D5A" => data <= "00110";
                when x"D5B" => data <= "00000";
                when x"D5C" => data <= "00110";
                when x"D5D" => data <= "00000";
                when x"D5E" => data <= "00001";
                when x"D5F" => data <= "00110";
                when x"D60" => data <= "11000";
                when x"D61" => data <= "00000";
                when x"D62" => data <= "00000";
                when x"D63" => data <= "00000";
                when x"D64" => data <= "00000";
                when x"D65" => data <= "00000";
                when x"D66" => data <= "00110";
                when x"D67" => data <= "00110";
                when x"D68" => data <= "00110";
                when x"D69" => data <= "00000";
                when x"D6A" => data <= "00110";
                when x"D6B" => data <= "00000";
                when x"D6C" => data <= "00000";
                when x"D6D" => data <= "00000";
                when x"D6E" => data <= "00101";
                when x"D6F" => data <= "00110";
                when x"D70" => data <= "00000";
                when x"D71" => data <= "11100";
                when x"D72" => data <= "10000";
                when x"D73" => data <= "00110";
                when x"D74" => data <= "00110";
                when x"D75" => data <= "00110";
                when x"D76" => data <= "00110";
                when x"D77" => data <= "00110";
                when x"D78" => data <= "00000";
                when x"D79" => data <= "00110";
                when x"D7A" => data <= "11010";
                when x"D7B" => data <= "00110";
                when x"D7C" => data <= "00110";
                when x"D7D" => data <= "00110";
                when x"D7E" => data <= "00110";
                when x"D7F" => data <= "00000";
                when x"D80" => data <= "00000";
                when x"D81" => data <= "00110";
                when x"D82" => data <= "00110";
                when x"D83" => data <= "00000";
                when x"D84" => data <= "00110";
                when x"D85" => data <= "00110";
                when x"D86" => data <= "11000";
                when x"D87" => data <= "01110";
                when x"D88" => data <= "11110";
                when x"D89" => data <= "00110";
                when x"D8A" => data <= "00000";
                when x"D8B" => data <= "00110";
                when x"D8C" => data <= "00000";
                when x"D8D" => data <= "00110";
                when x"D8E" => data <= "01001";
                when x"D8F" => data <= "00110";
                when x"D90" => data <= "00000";
                when x"D91" => data <= "00110";
                when x"D92" => data <= "00000";
                when x"D93" => data <= "00000";
                when x"D94" => data <= "00110";
                when x"D95" => data <= "00000";
                when x"D96" => data <= "00000";
                when x"D97" => data <= "00000";
                when x"D98" => data <= "00110";
                when x"D99" => data <= "00110";
                when x"D9A" => data <= "00110";
                when x"D9B" => data <= "00110";
                when x"D9C" => data <= "00000";
                when x"D9D" => data <= "10101";
                when x"D9E" => data <= "11111";
                when x"D9F" => data <= "00110";
                when x"DA0" => data <= "00000";
                when x"DA1" => data <= "00110";
                when x"DA2" => data <= "00110";
                when x"DA3" => data <= "00000";
                when x"DA4" => data <= "00000";
                when x"DA5" => data <= "00110";
                when x"DA6" => data <= "00000";
                when x"DA7" => data <= "00000";
                when x"DA8" => data <= "00110";
                when x"DA9" => data <= "00000";
                when x"DAA" => data <= "00000";
                when x"DAB" => data <= "00110";
                when x"DAC" => data <= "00110";
                when x"DAD" => data <= "00110";
                when x"DAE" => data <= "00110";
                when x"DAF" => data <= "11000";
                when x"DB0" => data <= "00000";
                when x"DB1" => data <= "00110";
                when x"DB2" => data <= "11101";
                when x"DB3" => data <= "00110";
                when x"DB4" => data <= "00000";
                when x"DB5" => data <= "10110";
                when x"DB6" => data <= "00000";
                when x"DB7" => data <= "00110";
                when x"DB8" => data <= "00110";
                when x"DB9" => data <= "00000";
                when x"DBA" => data <= "00110";
                when x"DBB" => data <= "01100";
                when x"DBC" => data <= "10001";
                when x"DBD" => data <= "00000";
                when x"DBE" => data <= "00110";
                when x"DBF" => data <= "00110";
                when x"DC0" => data <= "01010";
                when x"DC1" => data <= "00000";
                when x"DC2" => data <= "00110";
                when x"DC3" => data <= "00000";
                when x"DC4" => data <= "01110";
                when x"DC5" => data <= "00000";
                when x"DC6" => data <= "00110";
                when x"DC7" => data <= "10111";
                when x"DC8" => data <= "00000";
                when x"DC9" => data <= "00110";
                when x"DCA" => data <= "00000";
                when x"DCB" => data <= "01110";
                when x"DCC" => data <= "00000";
                when x"DCD" => data <= "00000";
                when x"DCE" => data <= "00110";
                when x"DCF" => data <= "00011";
                when x"DD0" => data <= "00110";
                when x"DD1" => data <= "00110";
                when x"DD2" => data <= "00000";
                when x"DD3" => data <= "00110";
                when x"DD4" => data <= "00110";
                when x"DD5" => data <= "00110";
                when x"DD6" => data <= "00110";
                when x"DD7" => data <= "00110";
                when x"DD8" => data <= "01101";
                when x"DD9" => data <= "00100";
                when x"DDA" => data <= "10010";
                when x"DDB" => data <= "00110";
                when x"DDC" => data <= "00110";
                when x"DDD" => data <= "00110";
                when x"DDE" => data <= "00000";
                when x"DDF" => data <= "00000";
                when x"DE0" => data <= "01110";
                when x"DE1" => data <= "00000";
                when x"DE2" => data <= "00110";
                when x"DE3" => data <= "00110";
                when x"DE4" => data <= "10110";
                when x"DE5" => data <= "00111";
                when x"DE6" => data <= "00110";
                when x"DE7" => data <= "00110";
                when x"DE8" => data <= "00000";
                when x"DE9" => data <= "00000";
                when x"DEA" => data <= "00110";
                when x"DEB" => data <= "00110";
                when x"DEC" => data <= "00000";
                when x"DED" => data <= "00110";
                when x"DEE" => data <= "10100";
                when x"DEF" => data <= "00110";
                when x"DF0" => data <= "00000";
                when x"DF1" => data <= "01011";
                when x"DF2" => data <= "00000";
                when x"DF3" => data <= "00000";
                when x"DF4" => data <= "00110";
                when x"DF5" => data <= "00110";
                when x"DF6" => data <= "00000";
                when x"DF7" => data <= "00000";
                when x"DF8" => data <= "00000";
                when x"DF9" => data <= "11111";
                when x"DFA" => data <= "00110";
                when x"DFB" => data <= "00101";
                when x"DFC" => data <= "00110";
                when x"DFD" => data <= "00110";
                when x"DFE" => data <= "00110";
                when x"DFF" => data <= "11101";
                when x"E00" => data <= "00110";
                when x"E01" => data <= "00000";
                when x"E02" => data <= "00110";
                when x"E03" => data <= "00000";
                when x"E04" => data <= "00000";
                when x"E05" => data <= "00000";
                when x"E06" => data <= "00000";
                when x"E07" => data <= "00000";
                when x"E08" => data <= "00000";
                when x"E09" => data <= "01101";
                when x"E0A" => data <= "00110";
                when x"E0B" => data <= "00110";
                when x"E0C" => data <= "00000";
                when x"E0D" => data <= "00000";
                when x"E0E" => data <= "00110";
                when x"E0F" => data <= "00110";
                when x"E10" => data <= "00000";
                when x"E11" => data <= "00011";
                when x"E12" => data <= "10101";
                when x"E13" => data <= "00110";
                when x"E14" => data <= "10011";
                when x"E15" => data <= "10011";
                when x"E16" => data <= "00000";
                when x"E17" => data <= "00000";
                when x"E18" => data <= "00000";
                when x"E19" => data <= "01000";
                when x"E1A" => data <= "00110";
                when x"E1B" => data <= "00100";
                when x"E1C" => data <= "00110";
                when x"E1D" => data <= "00000";
                when x"E1E" => data <= "01010";
                when x"E1F" => data <= "00000";
                when x"E20" => data <= "01000";
                when x"E21" => data <= "00000";
                when x"E22" => data <= "00110";
                when x"E23" => data <= "00110";
                when x"E24" => data <= "01000";
                when x"E25" => data <= "00110";
                when x"E26" => data <= "00000";
                when x"E27" => data <= "00110";
                when x"E28" => data <= "00000";
                when x"E29" => data <= "00110";
                when x"E2A" => data <= "00110";
                when x"E2B" => data <= "00110";
                when x"E2C" => data <= "00110";
                when x"E2D" => data <= "00000";
                when x"E2E" => data <= "00110";
                when x"E2F" => data <= "00000";
                when x"E30" => data <= "00000";
                when x"E31" => data <= "00110";
                when x"E32" => data <= "00000";
                when x"E33" => data <= "00000";
                when x"E34" => data <= "00110";
                when x"E35" => data <= "00110";
                when x"E36" => data <= "00000";
                when x"E37" => data <= "00000";
                when x"E38" => data <= "00000";
                when x"E39" => data <= "01101";
                when x"E3A" => data <= "00110";
                when x"E3B" => data <= "00110";
                when x"E3C" => data <= "00110";
                when x"E3D" => data <= "00110";
                when x"E3E" => data <= "00001";
                when x"E3F" => data <= "00011";
                when x"E40" => data <= "00000";
                when x"E41" => data <= "00000";
                when x"E42" => data <= "00110";
                when x"E43" => data <= "00000";
                when x"E44" => data <= "00011";
                when x"E45" => data <= "11011";
                when x"E46" => data <= "11001";
                when x"E47" => data <= "10011";
                when x"E48" => data <= "00110";
                when x"E49" => data <= "00000";
                when x"E4A" => data <= "00110";
                when x"E4B" => data <= "00110";
                when x"E4C" => data <= "00000";
                when x"E4D" => data <= "00000";
                when x"E4E" => data <= "00010";
                when x"E4F" => data <= "00110";
                when x"E50" => data <= "00000";
                when x"E51" => data <= "00110";
                when x"E52" => data <= "00110";
                when x"E53" => data <= "00110";
                when x"E54" => data <= "10111";
                when x"E55" => data <= "00110";
                when x"E56" => data <= "00000";
                when x"E57" => data <= "00000";
                when x"E58" => data <= "00000";
                when x"E59" => data <= "01011";
                when x"E5A" => data <= "00000";
                when x"E5B" => data <= "11000";
                when x"E5C" => data <= "00000";
                when x"E5D" => data <= "00000";
                when x"E5E" => data <= "00000";
                when x"E5F" => data <= "00110";
                when x"E60" => data <= "00110";
                when x"E61" => data <= "00110";
                when x"E62" => data <= "00110";
                when x"E63" => data <= "00110";
                when x"E64" => data <= "00000";
                when x"E65" => data <= "00110";
                when x"E66" => data <= "00000";
                when x"E67" => data <= "00110";
                when x"E68" => data <= "00110";
                when x"E69" => data <= "00110";
                when x"E6A" => data <= "00110";
                when x"E6B" => data <= "00011";
                when x"E6C" => data <= "00000";
                when x"E6D" => data <= "11001";
                when x"E6E" => data <= "00000";
                when x"E6F" => data <= "00000";
                when x"E70" => data <= "00110";
                when x"E71" => data <= "00000";
                when x"E72" => data <= "10111";
                when x"E73" => data <= "00000";
                when x"E74" => data <= "00000";
                when x"E75" => data <= "00000";
                when x"E76" => data <= "00000";
                when x"E77" => data <= "00110";
                when x"E78" => data <= "00110";
                when x"E79" => data <= "11001";
                when x"E7A" => data <= "00000";
                when x"E7B" => data <= "00000";
                when x"E7C" => data <= "00000";
                when x"E7D" => data <= "01011";
                when x"E7E" => data <= "00000";
                when x"E7F" => data <= "00110";
                when x"E80" => data <= "00000";
                when x"E81" => data <= "00110";
                when x"E82" => data <= "00000";
                when x"E83" => data <= "00110";
                when x"E84" => data <= "00110";
                when x"E85" => data <= "00000";
                when x"E86" => data <= "00000";
                when x"E87" => data <= "00110";
                when x"E88" => data <= "00010";
                when x"E89" => data <= "00110";
                when x"E8A" => data <= "00110";
                when x"E8B" => data <= "00000";
                when x"E8C" => data <= "00000";
                when x"E8D" => data <= "00000";
                when x"E8E" => data <= "01010";
                when x"E8F" => data <= "00110";
                when x"E90" => data <= "00110";
                when x"E91" => data <= "01111";
                when x"E92" => data <= "11110";
                when x"E93" => data <= "00111";
                when x"E94" => data <= "00000";
                when x"E95" => data <= "00110";
                when x"E96" => data <= "00000";
                when x"E97" => data <= "00110";
                when x"E98" => data <= "00111";
                when x"E99" => data <= "00000";
                when x"E9A" => data <= "00110";
                when x"E9B" => data <= "00000";
                when x"E9C" => data <= "00000";
                when x"E9D" => data <= "00110";
                when x"E9E" => data <= "00000";
                when x"E9F" => data <= "00110";
                when x"EA0" => data <= "00000";
                when x"EA1" => data <= "10010";
                when x"EA2" => data <= "00000";
                when x"EA3" => data <= "00110";
                when x"EA4" => data <= "00110";
                when x"EA5" => data <= "00101";
                when x"EA6" => data <= "00000";
                when x"EA7" => data <= "00000";
                when x"EA8" => data <= "00110";
                when x"EA9" => data <= "00011";
                when x"EAA" => data <= "00110";
                when x"EAB" => data <= "00000";
                when x"EAC" => data <= "00000";
                when x"EAD" => data <= "01101";
                when x"EAE" => data <= "00100";
                when x"EAF" => data <= "00000";
                when x"EB0" => data <= "01101";
                when x"EB1" => data <= "00000";
                when x"EB2" => data <= "10101";
                when x"EB3" => data <= "00110";
                when x"EB4" => data <= "00110";
                when x"EB5" => data <= "00000";
                when x"EB6" => data <= "00110";
                when x"EB7" => data <= "00110";
                when x"EB8" => data <= "00000";
                when x"EB9" => data <= "00110";
                when x"EBA" => data <= "00110";
                when x"EBB" => data <= "10101";
                when x"EBC" => data <= "00000";
                when x"EBD" => data <= "00110";
                when x"EBE" => data <= "01101";
                when x"EBF" => data <= "00000";
                when x"EC0" => data <= "00000";
                when x"EC1" => data <= "01101";
                when x"EC2" => data <= "00110";
                when x"EC3" => data <= "00110";
                when x"EC4" => data <= "00110";
                when x"EC5" => data <= "00000";
                when x"EC6" => data <= "00000";
                when x"EC7" => data <= "00000";
                when x"EC8" => data <= "00110";
                when x"EC9" => data <= "00110";
                when x"ECA" => data <= "00110";
                when x"ECB" => data <= "10101";
                when x"ECC" => data <= "01110";
                when x"ECD" => data <= "00000";
                when x"ECE" => data <= "00000";
                when x"ECF" => data <= "00110";
                when x"ED0" => data <= "11100";
                when x"ED1" => data <= "00000";
                when x"ED2" => data <= "00000";
                when x"ED3" => data <= "00110";
                when x"ED4" => data <= "00110";
                when x"ED5" => data <= "00110";
                when x"ED6" => data <= "00000";
                when x"ED7" => data <= "01001";
                when x"ED8" => data <= "00110";
                when x"ED9" => data <= "00000";
                when x"EDA" => data <= "00110";
                when x"EDB" => data <= "00000";
                when x"EDC" => data <= "00110";
                when x"EDD" => data <= "00000";
                when x"EDE" => data <= "00000";
                when x"EDF" => data <= "10101";
                when x"EE0" => data <= "00000";
                when x"EE1" => data <= "00000";
                when x"EE2" => data <= "00000";
                when x"EE3" => data <= "01100";
                when x"EE4" => data <= "00110";
                when x"EE5" => data <= "01101";
                when x"EE6" => data <= "10001";
                when x"EE7" => data <= "00110";
                when x"EE8" => data <= "10111";
                when x"EE9" => data <= "00110";
                when x"EEA" => data <= "00111";
                when x"EEB" => data <= "00000";
                when x"EEC" => data <= "11100";
                when x"EED" => data <= "00000";
                when x"EEE" => data <= "00110";
                when x"EEF" => data <= "00110";
                when x"EF0" => data <= "00000";
                when x"EF1" => data <= "00110";
                when x"EF2" => data <= "10111";
                when x"EF3" => data <= "00110";
                when x"EF4" => data <= "00110";
                when x"EF5" => data <= "00000";
                when x"EF6" => data <= "10001";
                when x"EF7" => data <= "00000";
                when x"EF8" => data <= "00110";
                when x"EF9" => data <= "00110";
                when x"EFA" => data <= "00110";
                when x"EFB" => data <= "00110";
                when x"EFC" => data <= "00110";
                when x"EFD" => data <= "00110";
                when x"EFE" => data <= "00110";
                when x"EFF" => data <= "00000";
                when x"F00" => data <= "00110";
                when x"F01" => data <= "00110";
                when x"F02" => data <= "00000";
                when x"F03" => data <= "00110";
                when x"F04" => data <= "00000";
                when x"F05" => data <= "00000";
                when x"F06" => data <= "00110";
                when x"F07" => data <= "00110";
                when x"F08" => data <= "00000";
                when x"F09" => data <= "00110";
                when x"F0A" => data <= "00000";
                when x"F0B" => data <= "00000";
                when x"F0C" => data <= "00000";
                when x"F0D" => data <= "00110";
                when x"F0E" => data <= "00110";
                when x"F0F" => data <= "00000";
                when x"F10" => data <= "00000";
                when x"F11" => data <= "00110";
                when x"F12" => data <= "00000";
                when x"F13" => data <= "00110";
                when x"F14" => data <= "00000";
                when x"F15" => data <= "00000";
                when x"F16" => data <= "00000";
                when x"F17" => data <= "00000";
                when x"F18" => data <= "00000";
                when x"F19" => data <= "00110";
                when x"F1A" => data <= "00110";
                when x"F1B" => data <= "00110";
                when x"F1C" => data <= "00000";
                when x"F1D" => data <= "00000";
                when x"F1E" => data <= "00110";
                when x"F1F" => data <= "00110";
                when x"F20" => data <= "00110";
                when x"F21" => data <= "01011";
                when x"F22" => data <= "00000";
                when x"F23" => data <= "00110";
                when x"F24" => data <= "00110";
                when x"F25" => data <= "00000";
                when x"F26" => data <= "11101";
                when x"F27" => data <= "00000";
                when x"F28" => data <= "00110";
                when x"F29" => data <= "00110";
                when x"F2A" => data <= "00110";
                when x"F2B" => data <= "00000";
                when x"F2C" => data <= "00000";
                when x"F2D" => data <= "11000";
                when x"F2E" => data <= "00110";
                when x"F2F" => data <= "00110";
                when x"F30" => data <= "00000";
                when x"F31" => data <= "00000";
                when x"F32" => data <= "01101";
                when x"F33" => data <= "00000";
                when x"F34" => data <= "00110";
                when x"F35" => data <= "11111";
                when x"F36" => data <= "00000";
                when x"F37" => data <= "00000";
                when x"F38" => data <= "00110";
                when x"F39" => data <= "00000";
                when x"F3A" => data <= "00110";
                when x"F3B" => data <= "00110";
                when x"F3C" => data <= "00110";
                when x"F3D" => data <= "01011";
                when x"F3E" => data <= "00000";
                when x"F3F" => data <= "00000";
                when x"F40" => data <= "00110";
                when x"F41" => data <= "00110";
                when x"F42" => data <= "00000";
                when x"F43" => data <= "00110";
                when x"F44" => data <= "00110";
                when x"F45" => data <= "00110";
                when x"F46" => data <= "00000";
                when x"F47" => data <= "00000";
                when x"F48" => data <= "00110";
                when x"F49" => data <= "00110";
                when x"F4A" => data <= "00110";
                when x"F4B" => data <= "11010";
                when x"F4C" => data <= "10111";
                when x"F4D" => data <= "00110";
                when x"F4E" => data <= "10000";
                when x"F4F" => data <= "00010";
                when x"F50" => data <= "00110";
                when x"F51" => data <= "00110";
                when x"F52" => data <= "00000";
                when x"F53" => data <= "00000";
                when x"F54" => data <= "00110";
                when x"F55" => data <= "10111";
                when x"F56" => data <= "01101";
                when x"F57" => data <= "00000";
                when x"F58" => data <= "11010";
                when x"F59" => data <= "00110";
                when x"F5A" => data <= "00000";
                when x"F5B" => data <= "00000";
                when x"F5C" => data <= "00000";
                when x"F5D" => data <= "00110";
                when x"F5E" => data <= "00000";
                when x"F5F" => data <= "00000";
                when x"F60" => data <= "00010";
                when x"F61" => data <= "01101";
                when x"F62" => data <= "11001";
                when x"F63" => data <= "00000";
                when x"F64" => data <= "00110";
                when x"F65" => data <= "00000";
                when x"F66" => data <= "00000";
                when x"F67" => data <= "00000";
                when x"F68" => data <= "10101";
                when x"F69" => data <= "00000";
                when x"F6A" => data <= "00110";
                when x"F6B" => data <= "10101";
                when x"F6C" => data <= "00110";
                when x"F6D" => data <= "10011";
                when x"F6E" => data <= "00110";
                when x"F6F" => data <= "00000";
                when x"F70" => data <= "00000";
                when x"F71" => data <= "00000";
                when x"F72" => data <= "00010";
                when x"F73" => data <= "00110";
                when x"F74" => data <= "00000";
                when x"F75" => data <= "00110";
                when x"F76" => data <= "00000";
                when x"F77" => data <= "00110";
                when x"F78" => data <= "00010";
                when x"F79" => data <= "00000";
                when x"F7A" => data <= "00000";
                when x"F7B" => data <= "10110";
                when x"F7C" => data <= "00000";
                when x"F7D" => data <= "00110";
                when x"F7E" => data <= "00000";
                when x"F7F" => data <= "00000";
                when x"F80" => data <= "00110";
                when x"F81" => data <= "00000";
                when x"F82" => data <= "01110";
                when x"F83" => data <= "00110";
                when x"F84" => data <= "10100";
                when x"F85" => data <= "00000";
                when x"F86" => data <= "00110";
                when x"F87" => data <= "00110";
                when x"F88" => data <= "00000";
                when x"F89" => data <= "01100";
                when x"F8A" => data <= "00000";
                when x"F8B" => data <= "00000";
                when x"F8C" => data <= "00110";
                when x"F8D" => data <= "00000";
                when x"F8E" => data <= "11101";
                when x"F8F" => data <= "00110";
                when x"F90" => data <= "00000";
                when x"F91" => data <= "00000";
                when x"F92" => data <= "00110";
                when x"F93" => data <= "11001";
                when x"F94" => data <= "01101";
                when x"F95" => data <= "00110";
                when x"F96" => data <= "00000";
                when x"F97" => data <= "00000";
                when x"F98" => data <= "10110";
                when x"F99" => data <= "00000";
                when x"F9A" => data <= "00110";
                when x"F9B" => data <= "11111";
                when x"F9C" => data <= "00000";
                when x"F9D" => data <= "10101";
                when x"F9E" => data <= "00110";
                when x"F9F" => data <= "00110";
                when x"FA0" => data <= "00000";
                when x"FA1" => data <= "00110";
                when x"FA2" => data <= "01011";
                when x"FA3" => data <= "00000";
                when x"FA4" => data <= "00000";
                when x"FA5" => data <= "00000";
                when x"FA6" => data <= "00000";
                when x"FA7" => data <= "01100";
                when x"FA8" => data <= "00110";
                when x"FA9" => data <= "10111";
                when x"FAA" => data <= "00000";
                when x"FAB" => data <= "00110";
                when x"FAC" => data <= "00000";
                when x"FAD" => data <= "00110";
                when x"FAE" => data <= "00000";
                when x"FAF" => data <= "00110";
                when x"FB0" => data <= "01011";
                when x"FB1" => data <= "00110";
                when x"FB2" => data <= "01010";
                when x"FB3" => data <= "00110";
                when x"FB4" => data <= "00110";
                when x"FB5" => data <= "00110";
                when x"FB6" => data <= "00000";
                when x"FB7" => data <= "10101";
                when x"FB8" => data <= "00000";
                when x"FB9" => data <= "01001";
                when x"FBA" => data <= "00110";
                when x"FBB" => data <= "00110";
                when x"FBC" => data <= "00000";
                when x"FBD" => data <= "00000";
                when x"FBE" => data <= "00110";
                when x"FBF" => data <= "10001";
                when x"FC0" => data <= "00110";
                when x"FC1" => data <= "00110";
                when x"FC2" => data <= "10011";
                when x"FC3" => data <= "00000";
                when x"FC4" => data <= "00110";
                when x"FC5" => data <= "00000";
                when x"FC6" => data <= "00110";
                when x"FC7" => data <= "10001";
                when x"FC8" => data <= "00110";
                when x"FC9" => data <= "11001";
                when x"FCA" => data <= "00000";
                when x"FCB" => data <= "00110";
                when x"FCC" => data <= "00010";
                when x"FCD" => data <= "11001";
                when x"FCE" => data <= "00000";
                when x"FCF" => data <= "00000";
                when x"FD0" => data <= "00010";
                when x"FD1" => data <= "00110";
                when x"FD2" => data <= "11111";
                when x"FD3" => data <= "00110";
                when x"FD4" => data <= "11010";
                when x"FD5" => data <= "10101";
                when x"FD6" => data <= "00110";
                when x"FD7" => data <= "00110";
                when x"FD8" => data <= "00000";
                when x"FD9" => data <= "00110";
                when x"FDA" => data <= "10101";
                when x"FDB" => data <= "00110";
                when x"FDC" => data <= "01101";
                when x"FDD" => data <= "00000";
                when x"FDE" => data <= "01101";
                when x"FDF" => data <= "00110";
                when x"FE0" => data <= "00110";
                when x"FE1" => data <= "00000";
                when x"FE2" => data <= "11001";
                when x"FE3" => data <= "00110";
                when x"FE4" => data <= "00110";
                when x"FE5" => data <= "00110";
                when x"FE6" => data <= "00000";
                when x"FE7" => data <= "00000";
                when x"FE8" => data <= "00110";
                when x"FE9" => data <= "00000";
                when x"FEA" => data <= "00000";
                when x"FEB" => data <= "00110";
                when x"FEC" => data <= "10010";
                when x"FED" => data <= "00110";
                when x"FEE" => data <= "00000";
                when x"FEF" => data <= "00110";
                when x"FF0" => data <= "00110";
                when x"FF1" => data <= "00000";
                when x"FF2" => data <= "00110";
                when x"FF3" => data <= "00110";
                when x"FF4" => data <= "11000";
                when x"FF5" => data <= "01101";
                when x"FF6" => data <= "00110";
                when x"FF7" => data <= "00110";
                when x"FF8" => data <= "00110";
                when x"FF9" => data <= "00000";
                when x"FFA" => data <= "10111";
                when x"FFB" => data <= "00110";
                when x"FFC" => data <= "00110";
                when x"FFD" => data <= "10010";
                when x"FFE" => data <= "00000";
                when x"FFF" => data <= "00110";
                when x"1000" => data <= "00000";
                when x"1001" => data <= "00000";
                when x"1002" => data <= "00000";
                when x"1003" => data <= "00000";
                when x"1004" => data <= "00110";
                when x"1005" => data <= "01001";
                when x"1006" => data <= "00110";
                when x"1007" => data <= "00000";
                when x"1008" => data <= "10111";
                when x"1009" => data <= "00110";
                when x"100A" => data <= "00000";
                when x"100B" => data <= "00110";
                when x"100C" => data <= "00110";
                when x"100D" => data <= "01110";
                when x"100E" => data <= "00000";
                when x"100F" => data <= "00000";
                when x"1010" => data <= "00000";
                when x"1011" => data <= "00000";
                when x"1012" => data <= "00110";
                when x"1013" => data <= "00110";
                when x"1014" => data <= "00000";
                when x"1015" => data <= "00110";
                when x"1016" => data <= "00000";
                when x"1017" => data <= "00000";
                when x"1018" => data <= "00110";
                when x"1019" => data <= "10110";
                when x"101A" => data <= "00000";
                when x"101B" => data <= "00110";
                when x"101C" => data <= "00000";
                when x"101D" => data <= "00000";
                when x"101E" => data <= "00000";
                when x"101F" => data <= "00110";
                when x"1020" => data <= "00110";
                when x"1021" => data <= "00000";
                when x"1022" => data <= "00000";
                when x"1023" => data <= "00000";
                when x"1024" => data <= "11100";
                when x"1025" => data <= "00110";
                when x"1026" => data <= "00000";
                when x"1027" => data <= "00000";
                when x"1028" => data <= "00000";
                when x"1029" => data <= "00110";
                when x"102A" => data <= "01100";
                when x"102B" => data <= "00000";
                when x"102C" => data <= "00000";
                when x"102D" => data <= "00000";
                when x"102E" => data <= "00000";
                when x"102F" => data <= "11110";
                when x"1030" => data <= "00110";
                when x"1031" => data <= "00110";
                when x"1032" => data <= "00000";
                when x"1033" => data <= "00110";
                when x"1034" => data <= "00000";
                when x"1035" => data <= "01101";
                when x"1036" => data <= "01101";
                when x"1037" => data <= "11110";
                when x"1038" => data <= "00110";
                when x"1039" => data <= "10101";
                when x"103A" => data <= "00110";
                when x"103B" => data <= "00110";
                when x"103C" => data <= "00110";
                when x"103D" => data <= "00110";
                when x"103E" => data <= "00110";
                when x"103F" => data <= "00000";
                when x"1040" => data <= "11110";
                when x"1041" => data <= "00000";
                when x"1042" => data <= "00110";
                when x"1043" => data <= "10000";
                when x"1044" => data <= "00110";
                when x"1045" => data <= "00000";
                when x"1046" => data <= "00000";
                when x"1047" => data <= "00110";
                when x"1048" => data <= "00110";
                when x"1049" => data <= "01101";
                when x"104A" => data <= "01010";
                when x"104B" => data <= "00000";
                when x"104C" => data <= "01101";
                when x"104D" => data <= "00000";
                when x"104E" => data <= "00000";
                when x"104F" => data <= "10011";
                when x"1050" => data <= "00110";
                when x"1051" => data <= "00110";
                when x"1052" => data <= "00110";
                when x"1053" => data <= "00110";
                when x"1054" => data <= "00110";
                when x"1055" => data <= "00000";
                when x"1056" => data <= "00000";
                when x"1057" => data <= "01001";
                when x"1058" => data <= "00000";
                when x"1059" => data <= "00000";
                when x"105A" => data <= "00000";
                when x"105B" => data <= "00110";
                when x"105C" => data <= "00000";
                when x"105D" => data <= "10101";
                when x"105E" => data <= "00000";
                when x"105F" => data <= "00110";
                when x"1060" => data <= "00110";
                when x"1061" => data <= "00000";
                when x"1062" => data <= "01101";
                when x"1063" => data <= "00110";
                when x"1064" => data <= "00110";
                when x"1065" => data <= "01011";
                when x"1066" => data <= "00110";
                when x"1067" => data <= "01110";
                when x"1068" => data <= "00110";
                when x"1069" => data <= "00110";
                when x"106A" => data <= "00110";
                when x"106B" => data <= "00111";
                when x"106C" => data <= "00000";
                when x"106D" => data <= "00110";
                when x"106E" => data <= "11001";
                when x"106F" => data <= "00000";
                when x"1070" => data <= "00110";
                when x"1071" => data <= "01010";
                when x"1072" => data <= "00000";
                when x"1073" => data <= "00110";
                when x"1074" => data <= "00000";
                when x"1075" => data <= "01100";
                when x"1076" => data <= "11000";
                when x"1077" => data <= "00110";
                when x"1078" => data <= "00000";
                when x"1079" => data <= "00110";
                when x"107A" => data <= "01100";
                when x"107B" => data <= "00000";
                when x"107C" => data <= "00000";
                when x"107D" => data <= "00110";
                when x"107E" => data <= "11111";
                when x"107F" => data <= "00000";
                when x"1080" => data <= "00000";
                when x"1081" => data <= "00110";
                when x"1082" => data <= "00110";
                when x"1083" => data <= "00110";
                when x"1084" => data <= "00110";
                when x"1085" => data <= "00110";
                when x"1086" => data <= "00000";
                when x"1087" => data <= "00110";
                when x"1088" => data <= "00000";
                when x"1089" => data <= "00000";
                when x"108A" => data <= "00000";
                when x"108B" => data <= "00110";
                when x"108C" => data <= "00000";
                when x"108D" => data <= "00000";
                when x"108E" => data <= "11111";
                when x"108F" => data <= "10111";
                when x"1090" => data <= "00000";
                when x"1091" => data <= "00000";
                when x"1092" => data <= "00110";
                when x"1093" => data <= "00110";
                when x"1094" => data <= "00000";
                when x"1095" => data <= "00000";
                when x"1096" => data <= "00000";
                when x"1097" => data <= "00110";
                when x"1098" => data <= "11111";
                when x"1099" => data <= "00000";
                when x"109A" => data <= "00110";
                when x"109B" => data <= "00000";
                when x"109C" => data <= "00000";
                when x"109D" => data <= "10001";
                when x"109E" => data <= "00000";
                when x"109F" => data <= "00110";
                when x"10A0" => data <= "00110";
                when x"10A1" => data <= "00001";
                when x"10A2" => data <= "11110";
                when x"10A3" => data <= "00110";
                when x"10A4" => data <= "00000";
                when x"10A5" => data <= "00110";
                when x"10A6" => data <= "11111";
                when x"10A7" => data <= "00110";
                when x"10A8" => data <= "00110";
                when x"10A9" => data <= "00111";
                when x"10AA" => data <= "11100";
                when x"10AB" => data <= "00000";
                when x"10AC" => data <= "01011";
                when x"10AD" => data <= "00110";
                when x"10AE" => data <= "00000";
                when x"10AF" => data <= "00000";
                when x"10B0" => data <= "00110";
                when x"10B1" => data <= "00110";
                when x"10B2" => data <= "00000";
                when x"10B3" => data <= "00110";
                when x"10B4" => data <= "00000";
                when x"10B5" => data <= "00000";
                when x"10B6" => data <= "00110";
                when x"10B7" => data <= "00000";
                when x"10B8" => data <= "11000";
                when x"10B9" => data <= "01101";
                when x"10BA" => data <= "00000";
                when x"10BB" => data <= "00000";
                when x"10BC" => data <= "00000";
                when x"10BD" => data <= "00110";
                when x"10BE" => data <= "00110";
                when x"10BF" => data <= "00010";
                when x"10C0" => data <= "00000";
                when x"10C1" => data <= "00000";
                when x"10C2" => data <= "01011";
                when x"10C3" => data <= "11111";
                when x"10C4" => data <= "10001";
                when x"10C5" => data <= "00110";
                when x"10C6" => data <= "00000";
                when x"10C7" => data <= "00110";
                when x"10C8" => data <= "00110";
                when x"10C9" => data <= "00000";
                when x"10CA" => data <= "00000";
                when x"10CB" => data <= "00110";
                when x"10CC" => data <= "00110";
                when x"10CD" => data <= "00110";
                when x"10CE" => data <= "00000";
                when x"10CF" => data <= "00110";
                when x"10D0" => data <= "00000";
                when x"10D1" => data <= "00000";
                when x"10D2" => data <= "00000";
                when x"10D3" => data <= "11000";
                when x"10D4" => data <= "00110";
                when x"10D5" => data <= "00000";
                when x"10D6" => data <= "00110";
                when x"10D7" => data <= "00110";
                when x"10D8" => data <= "00010";
                when x"10D9" => data <= "01011";
                when x"10DA" => data <= "00110";
                when x"10DB" => data <= "00110";
                when x"10DC" => data <= "00110";
                when x"10DD" => data <= "00000";
                when x"10DE" => data <= "00110";
                when x"10DF" => data <= "00110";
                when x"10E0" => data <= "01011";
                when x"10E1" => data <= "00110";
                when x"10E2" => data <= "01011";
                when x"10E3" => data <= "11111";
                when x"10E4" => data <= "00110";
                when x"10E5" => data <= "01110";
                when x"10E6" => data <= "10011";
                when x"10E7" => data <= "10001";
                when x"10E8" => data <= "01011";
                when x"10E9" => data <= "00000";
                when x"10EA" => data <= "00000";
                when x"10EB" => data <= "00110";
                when x"10EC" => data <= "00000";
                when x"10ED" => data <= "00110";
                when x"10EE" => data <= "00110";
                when x"10EF" => data <= "00110";
                when x"10F0" => data <= "00110";
                when x"10F1" => data <= "00000";
                when x"10F2" => data <= "00110";
                when x"10F3" => data <= "00000";
                when x"10F4" => data <= "00000";
                when x"10F5" => data <= "00110";
                when x"10F6" => data <= "00000";
                when x"10F7" => data <= "11010";
                when x"10F8" => data <= "00110";
                when x"10F9" => data <= "00000";
                when x"10FA" => data <= "00000";
                when x"10FB" => data <= "01010";
                when x"10FC" => data <= "00110";
                when x"10FD" => data <= "00110";
                when x"10FE" => data <= "00000";
                when x"10FF" => data <= "00110";
                when x"1100" => data <= "01100";
                when x"1101" => data <= "00110";
                when x"1102" => data <= "00000";
                when x"1103" => data <= "01010";
                when x"1104" => data <= "00110";
                when x"1105" => data <= "10110";
                when x"1106" => data <= "00000";
                when x"1107" => data <= "00000";
                when x"1108" => data <= "00000";
                when x"1109" => data <= "00101";
                when x"110A" => data <= "00110";
                when x"110B" => data <= "00000";
                when x"110C" => data <= "10000";
                when x"110D" => data <= "01010";
                when x"110E" => data <= "01011";
                when x"110F" => data <= "11001";
                when x"1110" => data <= "00000";
                when x"1111" => data <= "00000";
                when x"1112" => data <= "00110";
                when x"1113" => data <= "11111";
                when x"1114" => data <= "00000";
                when x"1115" => data <= "00110";
                when x"1116" => data <= "00110";
                when x"1117" => data <= "00000";
                when x"1118" => data <= "01001";
                when x"1119" => data <= "00000";
                when x"111A" => data <= "00110";
                when x"111B" => data <= "00000";
                when x"111C" => data <= "00000";
                when x"111D" => data <= "00110";
                when x"111E" => data <= "11101";
                when x"111F" => data <= "00000";
                when x"1120" => data <= "00000";
                when x"1121" => data <= "00000";
                when x"1122" => data <= "00110";
                when x"1123" => data <= "01110";
                when x"1124" => data <= "00011";
                when x"1125" => data <= "00110";
                when x"1126" => data <= "01011";
                when x"1127" => data <= "00000";
                when x"1128" => data <= "10001";
                when x"1129" => data <= "00100";
                when x"112A" => data <= "00110";
                when x"112B" => data <= "00110";
                when x"112C" => data <= "00110";
                when x"112D" => data <= "00110";
                when x"112E" => data <= "00110";
                when x"112F" => data <= "00110";
                when x"1130" => data <= "00110";
                when x"1131" => data <= "00110";
                when x"1132" => data <= "00000";
                when x"1133" => data <= "00110";
                when x"1134" => data <= "11101";
                when x"1135" => data <= "00110";
                when x"1136" => data <= "00000";
                when x"1137" => data <= "10101";
                when x"1138" => data <= "01100";
                when x"1139" => data <= "00001";
                when x"113A" => data <= "00110";
                when x"113B" => data <= "00110";
                when x"113C" => data <= "00000";
                when x"113D" => data <= "00110";
                when x"113E" => data <= "00110";
                when x"113F" => data <= "00110";
                when x"1140" => data <= "00000";
                when x"1141" => data <= "00000";
                when x"1142" => data <= "00000";
                when x"1143" => data <= "00110";
                when x"1144" => data <= "00000";
                when x"1145" => data <= "00110";
                when x"1146" => data <= "00000";
                when x"1147" => data <= "00110";
                when x"1148" => data <= "01001";
                when x"1149" => data <= "00000";
                when x"114A" => data <= "00000";
                when x"114B" => data <= "00110";
                when x"114C" => data <= "11010";
                when x"114D" => data <= "00000";
                when x"114E" => data <= "00110";
                when x"114F" => data <= "01011";
                when x"1150" => data <= "00110";
                when x"1151" => data <= "00110";
                when x"1152" => data <= "10001";
                when x"1153" => data <= "00000";
                when x"1154" => data <= "00110";
                when x"1155" => data <= "00110";
                when x"1156" => data <= "00110";
                when x"1157" => data <= "00000";
                when x"1158" => data <= "00110";
                when x"1159" => data <= "00110";
                when x"115A" => data <= "00000";
                when x"115B" => data <= "00110";
                when x"115C" => data <= "11001";
                when x"115D" => data <= "00110";
                when x"115E" => data <= "00000";
                when x"115F" => data <= "00000";
                when x"1160" => data <= "00000";
                when x"1161" => data <= "10001";
                when x"1162" => data <= "01001";
                when x"1163" => data <= "11010";
                when x"1164" => data <= "00110";
                when x"1165" => data <= "00000";
                when x"1166" => data <= "00000";
                when x"1167" => data <= "00110";
                when x"1168" => data <= "00000";
                when x"1169" => data <= "00000";
                when x"116A" => data <= "00000";
                when x"116B" => data <= "00000";
                when x"116C" => data <= "00110";
                when x"116D" => data <= "00000";
                when x"116E" => data <= "10110";
                when x"116F" => data <= "01000";
                when x"1170" => data <= "00110";
                when x"1171" => data <= "00110";
                when x"1172" => data <= "00110";
                when x"1173" => data <= "00000";
                when x"1174" => data <= "00000";
                when x"1175" => data <= "00110";
                when x"1176" => data <= "00110";
                when x"1177" => data <= "00111";
                when x"1178" => data <= "00110";
                when x"1179" => data <= "00000";
                when x"117A" => data <= "00000";
                when x"117B" => data <= "00000";
                when x"117C" => data <= "00110";
                when x"117D" => data <= "00110";
                when x"117E" => data <= "00000";
                when x"117F" => data <= "00000";
                when x"1180" => data <= "00000";
                when x"1181" => data <= "00110";
                when x"1182" => data <= "00110";
                when x"1183" => data <= "00000";
                when x"1184" => data <= "00000";
                when x"1185" => data <= "00000";
                when x"1186" => data <= "01101";
                when x"1187" => data <= "00110";
                when x"1188" => data <= "01011";
                when x"1189" => data <= "00011";
                when x"118A" => data <= "00110";
                when x"118B" => data <= "10100";
                when x"118C" => data <= "00110";
                when x"118D" => data <= "01101";
                when x"118E" => data <= "00110";
                when x"118F" => data <= "00000";
                when x"1190" => data <= "00000";
                when x"1191" => data <= "00000";
                when x"1192" => data <= "00111";
                when x"1193" => data <= "00000";
                when x"1194" => data <= "00000";
                when x"1195" => data <= "00000";
                when x"1196" => data <= "01101";
                when x"1197" => data <= "00000";
                when x"1198" => data <= "00110";
                when x"1199" => data <= "00000";
                when x"119A" => data <= "01101";
                when x"119B" => data <= "00110";
                when x"119C" => data <= "00000";
                when x"119D" => data <= "00110";
                when x"119E" => data <= "00000";
                when x"119F" => data <= "00011";
                when x"11A0" => data <= "00110";
                when x"11A1" => data <= "00000";
                when x"11A2" => data <= "01001";
                when x"11A3" => data <= "00110";
                when x"11A4" => data <= "00000";
                when x"11A5" => data <= "00110";
                when x"11A6" => data <= "00000";
                when x"11A7" => data <= "00001";
                when x"11A8" => data <= "00110";
                when x"11A9" => data <= "00110";
                when x"11AA" => data <= "00000";
                when x"11AB" => data <= "00010";
                when x"11AC" => data <= "00000";
                when x"11AD" => data <= "11111";
                when x"11AE" => data <= "00110";
                when x"11AF" => data <= "01110";
                when x"11B0" => data <= "00000";
                when x"11B1" => data <= "00000";
                when x"11B2" => data <= "00110";
                when x"11B3" => data <= "00110";
                when x"11B4" => data <= "00000";
                when x"11B5" => data <= "00111";
                when x"11B6" => data <= "00000";
                when x"11B7" => data <= "00000";
                when x"11B8" => data <= "00110";
                when x"11B9" => data <= "00110";
                when x"11BA" => data <= "00000";
                when x"11BB" => data <= "00000";
                when x"11BC" => data <= "00101";
                when x"11BD" => data <= "00000";
                when x"11BE" => data <= "00110";
                when x"11BF" => data <= "00000";
                when x"11C0" => data <= "01101";
                when x"11C1" => data <= "00000";
                when x"11C2" => data <= "00110";
                when x"11C3" => data <= "00111";
                when x"11C4" => data <= "00111";
                when x"11C5" => data <= "01001";
                when x"11C6" => data <= "00111";
                when x"11C7" => data <= "00000";
                when x"11C8" => data <= "11010";
                when x"11C9" => data <= "00110";
                when x"11CA" => data <= "00000";
                when x"11CB" => data <= "11111";
                when x"11CC" => data <= "00110";
                when x"11CD" => data <= "00111";
                when x"11CE" => data <= "00000";
                when x"11CF" => data <= "00110";
                when x"11D0" => data <= "00000";
                when x"11D1" => data <= "00011";
                when x"11D2" => data <= "00110";
                when x"11D3" => data <= "01011";
                when x"11D4" => data <= "00000";
                when x"11D5" => data <= "00000";
                when x"11D6" => data <= "00001";
                when x"11D7" => data <= "00000";
                when x"11D8" => data <= "00000";
                when x"11D9" => data <= "00000";
                when x"11DA" => data <= "00000";
                when x"11DB" => data <= "00000";
                when x"11DC" => data <= "01101";
                when x"11DD" => data <= "00000";
                when x"11DE" => data <= "00110";
                when x"11DF" => data <= "00000";
                when x"11E0" => data <= "00000";
                when x"11E1" => data <= "10111";
                when x"11E2" => data <= "00110";
                when x"11E3" => data <= "00000";
                when x"11E4" => data <= "00110";
                when x"11E5" => data <= "00110";
                when x"11E6" => data <= "00000";
                when x"11E7" => data <= "00110";
                when x"11E8" => data <= "00000";
                when x"11E9" => data <= "00110";
                when x"11EA" => data <= "00000";
                when x"11EB" => data <= "01111";
                when x"11EC" => data <= "10000";
                when x"11ED" => data <= "00000";
                when x"11EE" => data <= "00011";
                when x"11EF" => data <= "01110";
                when x"11F0" => data <= "11100";
                when x"11F1" => data <= "01101";
                when x"11F2" => data <= "00000";
                when x"11F3" => data <= "00110";
                when x"11F4" => data <= "00000";
                when x"11F5" => data <= "00110";
                when x"11F6" => data <= "00110";
                when x"11F7" => data <= "00000";
                when x"11F8" => data <= "00110";
                when x"11F9" => data <= "00110";
                when x"11FA" => data <= "00110";
                when x"11FB" => data <= "01101";
                when x"11FC" => data <= "01010";
                when x"11FD" => data <= "00010";
                when x"11FE" => data <= "01001";
                when x"11FF" => data <= "00000";
                when x"1200" => data <= "00000";
                when x"1201" => data <= "00000";
                when x"1202" => data <= "00110";
                when x"1203" => data <= "11001";
                when x"1204" => data <= "00000";
                when x"1205" => data <= "00000";
                when x"1206" => data <= "00110";
                when x"1207" => data <= "00110";
                when x"1208" => data <= "00000";
                when x"1209" => data <= "00110";
                when x"120A" => data <= "00110";
                when x"120B" => data <= "00110";
                when x"120C" => data <= "00110";
                when x"120D" => data <= "11011";
                when x"120E" => data <= "00000";
                when x"120F" => data <= "00000";
                when x"1210" => data <= "00000";
                when x"1211" => data <= "00000";
                when x"1212" => data <= "00000";
                when x"1213" => data <= "10101";
                when x"1214" => data <= "00000";
                when x"1215" => data <= "11010";
                when x"1216" => data <= "00110";
                when x"1217" => data <= "00110";
                when x"1218" => data <= "00110";
                when x"1219" => data <= "00110";
                when x"121A" => data <= "01010";
                when x"121B" => data <= "00000";
                when x"121C" => data <= "00110";
                when x"121D" => data <= "00000";
                when x"121E" => data <= "00000";
                when x"121F" => data <= "00110";
                when x"1220" => data <= "00110";
                when x"1221" => data <= "00000";
                when x"1222" => data <= "10101";
                when x"1223" => data <= "00110";
                when x"1224" => data <= "00000";
                when x"1225" => data <= "00000";
                when x"1226" => data <= "00000";
                when x"1227" => data <= "00010";
                when x"1228" => data <= "01010";
                when x"1229" => data <= "00000";
                when x"122A" => data <= "00110";
                when x"122B" => data <= "00000";
                when x"122C" => data <= "00110";
                when x"122D" => data <= "00000";
                when x"122E" => data <= "00000";
                when x"122F" => data <= "00110";
                when x"1230" => data <= "00000";
                when x"1231" => data <= "00000";
                when x"1232" => data <= "00110";
                when x"1233" => data <= "00000";
                when x"1234" => data <= "00000";
                when x"1235" => data <= "00110";
                when x"1236" => data <= "00110";
                when x"1237" => data <= "00000";
                when x"1238" => data <= "00110";
                when x"1239" => data <= "00000";
                when x"123A" => data <= "00110";
                when x"123B" => data <= "00110";
                when x"123C" => data <= "00110";
                when x"123D" => data <= "11001";
                when x"123E" => data <= "10101";
                when x"123F" => data <= "10011";
                when x"1240" => data <= "00000";
                when x"1241" => data <= "11111";
                when x"1242" => data <= "00000";
                when x"1243" => data <= "00000";
                when x"1244" => data <= "00110";
                when x"1245" => data <= "00000";
                when x"1246" => data <= "00110";
                when x"1247" => data <= "10011";
                when x"1248" => data <= "00110";
                when x"1249" => data <= "00110";
                when x"124A" => data <= "00110";
                when x"124B" => data <= "01111";
                when x"124C" => data <= "00110";
                when x"124D" => data <= "00110";
                when x"124E" => data <= "00000";
                when x"124F" => data <= "00110";
                when x"1250" => data <= "00110";
                when x"1251" => data <= "00000";
                when x"1252" => data <= "00110";
                when x"1253" => data <= "00101";
                when x"1254" => data <= "00110";
                when x"1255" => data <= "00110";
                when x"1256" => data <= "00000";
                when x"1257" => data <= "00110";
                when x"1258" => data <= "00000";
                when x"1259" => data <= "00000";
                when x"125A" => data <= "00000";
                when x"125B" => data <= "00110";
                when x"125C" => data <= "00110";
                when x"125D" => data <= "11110";
                when x"125E" => data <= "00000";
                when x"125F" => data <= "00110";
                when x"1260" => data <= "00000";
                when x"1261" => data <= "00000";
                when x"1262" => data <= "00110";
                when x"1263" => data <= "01111";
                when x"1264" => data <= "00110";
                when x"1265" => data <= "00110";
                when x"1266" => data <= "00000";
                when x"1267" => data <= "00000";
                when x"1268" => data <= "00000";
                when x"1269" => data <= "00000";
                when x"126A" => data <= "00110";
                when x"126B" => data <= "00000";
                when x"126C" => data <= "00000";
                when x"126D" => data <= "10011";
                when x"126E" => data <= "00000";
                when x"126F" => data <= "00000";
                when x"1270" => data <= "00000";
                when x"1271" => data <= "10111";
                when x"1272" => data <= "00110";
                when x"1273" => data <= "00000";
                when x"1274" => data <= "00000";
                when x"1275" => data <= "00000";
                when x"1276" => data <= "00000";
                when x"1277" => data <= "00110";
                when x"1278" => data <= "00110";
                when x"1279" => data <= "00110";
                when x"127A" => data <= "11010";
                when x"127B" => data <= "00000";
                when x"127C" => data <= "00000";
                when x"127D" => data <= "00110";
                when x"127E" => data <= "00110";
                when x"127F" => data <= "00110";
                when x"1280" => data <= "00110";
                when x"1281" => data <= "00110";
                when x"1282" => data <= "00110";
                when x"1283" => data <= "00000";
                when x"1284" => data <= "00110";
                when x"1285" => data <= "00000";
                when x"1286" => data <= "01000";
                when x"1287" => data <= "01101";
                when x"1288" => data <= "00000";
                when x"1289" => data <= "00000";
                when x"128A" => data <= "00000";
                when x"128B" => data <= "00000";
                when x"128C" => data <= "10010";
                when x"128D" => data <= "11111";
                when x"128E" => data <= "00000";
                when x"128F" => data <= "00000";
                when x"1290" => data <= "00110";
                when x"1291" => data <= "00110";
                when x"1292" => data <= "00000";
                when x"1293" => data <= "00000";
                when x"1294" => data <= "00000";
                when x"1295" => data <= "00110";
                when x"1296" => data <= "00000";
                when x"1297" => data <= "00110";
                when x"1298" => data <= "00000";
                when x"1299" => data <= "00000";
                when x"129A" => data <= "00110";
                when x"129B" => data <= "00000";
                when x"129C" => data <= "00110";
                when x"129D" => data <= "00000";
                when x"129E" => data <= "11001";
                when x"129F" => data <= "00110";
                when x"12A0" => data <= "00000";
                when x"12A1" => data <= "00000";
                when x"12A2" => data <= "00110";
                when x"12A3" => data <= "00000";
                when x"12A4" => data <= "00110";
                when x"12A5" => data <= "00000";
                when x"12A6" => data <= "00110";
                when x"12A7" => data <= "00000";
                when x"12A8" => data <= "00110";
                when x"12A9" => data <= "00000";
                when x"12AA" => data <= "00110";
                when x"12AB" => data <= "00110";
                when x"12AC" => data <= "00000";
                when x"12AD" => data <= "00110";
                when x"12AE" => data <= "00000";
                when x"12AF" => data <= "00000";
                when x"12B0" => data <= "00110";
                when x"12B1" => data <= "00000";
                when x"12B2" => data <= "01101";
                when x"12B3" => data <= "01011";
                when x"12B4" => data <= "00110";
                when x"12B5" => data <= "00110";
                when x"12B6" => data <= "01100";
                when x"12B7" => data <= "10000";
                when x"12B8" => data <= "00110";
                when x"12B9" => data <= "00000";
                when x"12BA" => data <= "00000";
                when x"12BB" => data <= "00110";
                when x"12BC" => data <= "00111";
                when x"12BD" => data <= "00110";
                when x"12BE" => data <= "00110";
                when x"12BF" => data <= "01100";
                when x"12C0" => data <= "00110";
                when x"12C1" => data <= "00000";
                when x"12C2" => data <= "11101";
                when x"12C3" => data <= "00111";
                when x"12C4" => data <= "00000";
                when x"12C5" => data <= "01100";
                when x"12C6" => data <= "11010";
                when x"12C7" => data <= "00110";
                when x"12C8" => data <= "00110";
                when x"12C9" => data <= "00000";
                when x"12CA" => data <= "00000";
                when x"12CB" => data <= "11111";
                when x"12CC" => data <= "00000";
                when x"12CD" => data <= "01111";
                when x"12CE" => data <= "00110";
                when x"12CF" => data <= "11010";
                when x"12D0" => data <= "00101";
                when x"12D1" => data <= "00000";
                when x"12D2" => data <= "00111";
                when x"12D3" => data <= "00110";
                when x"12D4" => data <= "00000";
                when x"12D5" => data <= "01011";
                when x"12D6" => data <= "00000";
                when x"12D7" => data <= "00000";
                when x"12D8" => data <= "00110";
                when x"12D9" => data <= "00010";
                when x"12DA" => data <= "00000";
                when x"12DB" => data <= "00000";
                when x"12DC" => data <= "00110";
                when x"12DD" => data <= "00000";
                when x"12DE" => data <= "01011";
                when x"12DF" => data <= "10110";
                when x"12E0" => data <= "00110";
                when x"12E1" => data <= "10101";
                when x"12E2" => data <= "01010";
                when x"12E3" => data <= "00000";
                when x"12E4" => data <= "00110";
                when x"12E5" => data <= "00110";
                when x"12E6" => data <= "00110";
                when x"12E7" => data <= "01011";
                when x"12E8" => data <= "00110";
                when x"12E9" => data <= "01110";
                when x"12EA" => data <= "00000";
                when x"12EB" => data <= "00110";
                when x"12EC" => data <= "00000";
                when x"12ED" => data <= "00000";
                when x"12EE" => data <= "00000";
                when x"12EF" => data <= "00110";
                when x"12F0" => data <= "11100";
                when x"12F1" => data <= "00110";
                when x"12F2" => data <= "01101";
                when x"12F3" => data <= "10101";
                when x"12F4" => data <= "01001";
                when x"12F5" => data <= "01000";
                when x"12F6" => data <= "00110";
                when x"12F7" => data <= "11110";
                when x"12F8" => data <= "00110";
                when x"12F9" => data <= "00000";
                when x"12FA" => data <= "00110";
                when x"12FB" => data <= "00000";
                when x"12FC" => data <= "10000";
                when x"12FD" => data <= "01001";
                when x"12FE" => data <= "00000";
                when x"12FF" => data <= "00110";
                when x"1300" => data <= "00000";
                when x"1301" => data <= "00000";
                when x"1302" => data <= "00000";
                when x"1303" => data <= "00000";
                when x"1304" => data <= "00011";
                when x"1305" => data <= "00110";
                when x"1306" => data <= "00110";
                when x"1307" => data <= "00000";
                when x"1308" => data <= "00110";
                when x"1309" => data <= "01001";
                when x"130A" => data <= "11000";
                when x"130B" => data <= "00000";
                when x"130C" => data <= "11101";
                when x"130D" => data <= "00110";
                when x"130E" => data <= "00110";
                when x"130F" => data <= "00000";
                when x"1310" => data <= "00110";
                when x"1311" => data <= "00110";
                when x"1312" => data <= "00110";
                when x"1313" => data <= "00000";
                when x"1314" => data <= "01101";
                when x"1315" => data <= "00110";
                when x"1316" => data <= "01010";
                when x"1317" => data <= "00000";
                when x"1318" => data <= "00110";
                when x"1319" => data <= "00110";
                when x"131A" => data <= "00000";
                when x"131B" => data <= "00000";
                when x"131C" => data <= "00000";
                when x"131D" => data <= "00000";
                when x"131E" => data <= "00110";
                when x"131F" => data <= "00000";
                when x"1320" => data <= "00000";
                when x"1321" => data <= "00111";
                when x"1322" => data <= "00110";
                when x"1323" => data <= "00110";
                when x"1324" => data <= "00000";
                when x"1325" => data <= "00000";
                when x"1326" => data <= "00000";
                when x"1327" => data <= "00110";
                when x"1328" => data <= "00000";
                when x"1329" => data <= "00101";
                when x"132A" => data <= "00110";
                when x"132B" => data <= "00000";
                when x"132C" => data <= "10100";
                when x"132D" => data <= "00000";
                when x"132E" => data <= "00110";
                when x"132F" => data <= "00000";
                when x"1330" => data <= "11100";
                when x"1331" => data <= "00110";
                when x"1332" => data <= "00001";
                when x"1333" => data <= "00000";
                when x"1334" => data <= "00000";
                when x"1335" => data <= "00001";
                when x"1336" => data <= "00000";
                when x"1337" => data <= "00010";
                when x"1338" => data <= "00110";
                when x"1339" => data <= "00000";
                when x"133A" => data <= "00000";
                when x"133B" => data <= "00000";
                when x"133C" => data <= "00000";
                when x"133D" => data <= "00110";
                when x"133E" => data <= "01011";
                when x"133F" => data <= "00000";
                when x"1340" => data <= "00011";
                when x"1341" => data <= "10011";
                when x"1342" => data <= "00110";
                when x"1343" => data <= "00000";
                when x"1344" => data <= "00000";
                when x"1345" => data <= "00000";
                when x"1346" => data <= "00000";
                when x"1347" => data <= "01101";
                when x"1348" => data <= "10100";
                when x"1349" => data <= "00110";
                when x"134A" => data <= "00000";
                when x"134B" => data <= "00000";
                when x"134C" => data <= "00110";
                when x"134D" => data <= "00000";
                when x"134E" => data <= "00110";
                when x"134F" => data <= "00110";
                when x"1350" => data <= "00000";
                when x"1351" => data <= "00000";
                when x"1352" => data <= "00000";
                when x"1353" => data <= "00000";
                when x"1354" => data <= "00110";
                when x"1355" => data <= "00000";
                when x"1356" => data <= "00110";
                when x"1357" => data <= "11010";
                when x"1358" => data <= "00110";
                when x"1359" => data <= "00000";
                when x"135A" => data <= "00110";
                when x"135B" => data <= "00110";
                when x"135C" => data <= "00000";
                when x"135D" => data <= "00110";
                when x"135E" => data <= "00000";
                when x"135F" => data <= "00000";
                when x"1360" => data <= "01010";
                when x"1361" => data <= "00110";
                when x"1362" => data <= "00000";
                when x"1363" => data <= "00110";
                when x"1364" => data <= "00110";
                when x"1365" => data <= "01110";
                when x"1366" => data <= "00110";
                when x"1367" => data <= "00110";
                when x"1368" => data <= "00000";
                when x"1369" => data <= "00110";
                when x"136A" => data <= "00000";
                when x"136B" => data <= "01101";
                when x"136C" => data <= "00110";
                when x"136D" => data <= "00110";
                when x"136E" => data <= "11111";
                when x"136F" => data <= "00000";
                when x"1370" => data <= "00000";
                when x"1371" => data <= "00000";
                when x"1372" => data <= "00110";
                when x"1373" => data <= "00110";
                when x"1374" => data <= "01010";
                when x"1375" => data <= "01011";
                when x"1376" => data <= "00111";
                when x"1377" => data <= "00000";
                when x"1378" => data <= "00110";
                when x"1379" => data <= "00110";
                when x"137A" => data <= "00110";
                when x"137B" => data <= "00000";
                when x"137C" => data <= "00000";
                when x"137D" => data <= "11001";
                when x"137E" => data <= "00000";
                when x"137F" => data <= "00110";
                when x"1380" => data <= "11010";
                when x"1381" => data <= "00000";
                when x"1382" => data <= "00111";
                when x"1383" => data <= "00110";
                when x"1384" => data <= "00110";
                when x"1385" => data <= "01111";
                when x"1386" => data <= "11001";
                when x"1387" => data <= "00000";
                when x"1388" => data <= "00110";
                when x"1389" => data <= "00000";
                when x"138A" => data <= "00110";
                when x"138B" => data <= "00110";
                when x"138C" => data <= "00110";
                when x"138D" => data <= "00110";
                when x"138E" => data <= "00110";
                when x"138F" => data <= "00000";
                when x"1390" => data <= "00110";
                when x"1391" => data <= "11111";
                when x"1392" => data <= "00110";
                when x"1393" => data <= "00110";
                when x"1394" => data <= "00110";
                when x"1395" => data <= "00000";
                when x"1396" => data <= "00000";
                when x"1397" => data <= "00000";
                when x"1398" => data <= "01010";
                when x"1399" => data <= "11001";
                when x"139A" => data <= "00110";
                when x"139B" => data <= "00110";
                when x"139C" => data <= "00000";
                when x"139D" => data <= "11011";
                when x"139E" => data <= "00110";
                when x"139F" => data <= "00000";
                when x"13A0" => data <= "00001";
                when x"13A1" => data <= "00110";
                when x"13A2" => data <= "11010";
                when x"13A3" => data <= "00000";
                when x"13A4" => data <= "00000";
                when x"13A5" => data <= "00110";
                when x"13A6" => data <= "00000";
                when x"13A7" => data <= "00000";
                when x"13A8" => data <= "00110";
                when x"13A9" => data <= "00000";
                when x"13AA" => data <= "00000";
                when x"13AB" => data <= "00000";
                when x"13AC" => data <= "00110";
                when x"13AD" => data <= "00110";
                when x"13AE" => data <= "00110";
                when x"13AF" => data <= "11110";
                when x"13B0" => data <= "00000";
                when x"13B1" => data <= "00000";
                when x"13B2" => data <= "00000";
                when x"13B3" => data <= "00110";
                when x"13B4" => data <= "11010";
                when x"13B5" => data <= "00110";
                when x"13B6" => data <= "00000";
                when x"13B7" => data <= "00110";
                when x"13B8" => data <= "00110";
                when x"13B9" => data <= "00000";
                when x"13BA" => data <= "00000";
                when x"13BB" => data <= "00000";
                when x"13BC" => data <= "00000";
                when x"13BD" => data <= "00100";
                when x"13BE" => data <= "00000";
                when x"13BF" => data <= "01011";
                when x"13C0" => data <= "00110";
                when x"13C1" => data <= "00110";
                when x"13C2" => data <= "10111";
                when x"13C3" => data <= "00110";
                when x"13C4" => data <= "00110";
                when x"13C5" => data <= "00110";
                when x"13C6" => data <= "00000";
                when x"13C7" => data <= "00110";
                when x"13C8" => data <= "00110";
                when x"13C9" => data <= "00110";
                when x"13CA" => data <= "00000";
                when x"13CB" => data <= "00000";
                when x"13CC" => data <= "00110";
                when x"13CD" => data <= "00000";
                when x"13CE" => data <= "00110";
                when x"13CF" => data <= "00110";
                when x"13D0" => data <= "00000";
                when x"13D1" => data <= "01010";
                when x"13D2" => data <= "00110";
                when x"13D3" => data <= "00110";
                when x"13D4" => data <= "00110";
                when x"13D5" => data <= "11000";
                when x"13D6" => data <= "00110";
                when x"13D7" => data <= "00110";
                when x"13D8" => data <= "00110";
                when x"13D9" => data <= "00110";
                when x"13DA" => data <= "00000";
                when x"13DB" => data <= "00101";
                when x"13DC" => data <= "00110";
                when x"13DD" => data <= "00110";
                when x"13DE" => data <= "01011";
                when x"13DF" => data <= "00000";
                when x"13E0" => data <= "10000";
                when x"13E1" => data <= "00000";
                when x"13E2" => data <= "00000";
                when x"13E3" => data <= "00000";
                when x"13E4" => data <= "00110";
                when x"13E5" => data <= "00000";
                when x"13E6" => data <= "00110";
                when x"13E7" => data <= "01010";
                when x"13E8" => data <= "00110";
                when x"13E9" => data <= "00000";
                when x"13EA" => data <= "00000";
                when x"13EB" => data <= "00110";
                when x"13EC" => data <= "00000";
                when x"13ED" => data <= "01010";
                when x"13EE" => data <= "00110";
                when x"13EF" => data <= "00110";
                when x"13F0" => data <= "00000";
                when x"13F1" => data <= "00110";
                when x"13F2" => data <= "00110";
                when x"13F3" => data <= "00110";
                when x"13F4" => data <= "00110";
                when x"13F5" => data <= "00000";
                when x"13F6" => data <= "00000";
                when x"13F7" => data <= "00000";
                when x"13F8" => data <= "00110";
                when x"13F9" => data <= "00110";
                when x"13FA" => data <= "00000";
                when x"13FB" => data <= "00110";
                when x"13FC" => data <= "00000";
                when x"13FD" => data <= "00000";
                when x"13FE" => data <= "00000";
                when x"13FF" => data <= "00110";
                when x"1400" => data <= "00110";
                when x"1401" => data <= "11011";
                when x"1402" => data <= "00110";
                when x"1403" => data <= "00000";
                when x"1404" => data <= "00110";
                when x"1405" => data <= "00110";
                when x"1406" => data <= "00110";
                when x"1407" => data <= "11001";
                when x"1408" => data <= "00110";
                when x"1409" => data <= "11001";
                when x"140A" => data <= "00110";
                when x"140B" => data <= "00000";
                when x"140C" => data <= "10010";
                when x"140D" => data <= "00000";
                when x"140E" => data <= "11101";
                when x"140F" => data <= "00000";
                when x"1410" => data <= "00110";
                when x"1411" => data <= "00110";
                when x"1412" => data <= "00110";
                when x"1413" => data <= "01000";
                when x"1414" => data <= "00110";
                when x"1415" => data <= "00000";
                when x"1416" => data <= "01111";
                when x"1417" => data <= "00000";
                when x"1418" => data <= "00000";
                when x"1419" => data <= "00000";
                when x"141A" => data <= "00000";
                when x"141B" => data <= "00110";
                when x"141C" => data <= "11110";
                when x"141D" => data <= "00000";
                when x"141E" => data <= "00110";
                when x"141F" => data <= "00000";
                when x"1420" => data <= "00000";
                when x"1421" => data <= "10101";
                when x"1422" => data <= "00000";
                when x"1423" => data <= "00000";
                when x"1424" => data <= "10011";
                when x"1425" => data <= "00000";
                when x"1426" => data <= "00000";
                when x"1427" => data <= "00000";
                when x"1428" => data <= "00000";
                when x"1429" => data <= "10111";
                when x"142A" => data <= "11000";
                when x"142B" => data <= "00110";
                when x"142C" => data <= "00110";
                when x"142D" => data <= "00010";
                when x"142E" => data <= "00110";
                when x"142F" => data <= "00110";
                when x"1430" => data <= "00000";
                when x"1431" => data <= "00000";
                when x"1432" => data <= "00110";
                when x"1433" => data <= "00000";
                when x"1434" => data <= "00110";
                when x"1435" => data <= "10010";
                when x"1436" => data <= "00000";
                when x"1437" => data <= "00111";
                when x"1438" => data <= "00000";
                when x"1439" => data <= "00001";
                when x"143A" => data <= "00110";
                when x"143B" => data <= "00000";
                when x"143C" => data <= "00000";
                when x"143D" => data <= "00000";
                when x"143E" => data <= "00000";
                when x"143F" => data <= "00110";
                when x"1440" => data <= "00000";
                when x"1441" => data <= "00101";
                when x"1442" => data <= "11100";
                when x"1443" => data <= "00000";
                when x"1444" => data <= "00110";
                when x"1445" => data <= "01010";
                when x"1446" => data <= "00000";
                when x"1447" => data <= "00110";
                when x"1448" => data <= "00110";
                when x"1449" => data <= "01101";
                when x"144A" => data <= "11110";
                when x"144B" => data <= "00000";
                when x"144C" => data <= "00000";
                when x"144D" => data <= "00110";
                when x"144E" => data <= "00110";
                when x"144F" => data <= "00000";
                when x"1450" => data <= "11001";
                when x"1451" => data <= "00000";
                when x"1452" => data <= "01101";
                when x"1453" => data <= "11111";
                when x"1454" => data <= "00110";
                when x"1455" => data <= "00000";
                when x"1456" => data <= "00000";
                when x"1457" => data <= "00000";
                when x"1458" => data <= "01000";
                when x"1459" => data <= "00111";
                when x"145A" => data <= "01000";
                when x"145B" => data <= "00000";
                when x"145C" => data <= "10101";
                when x"145D" => data <= "01011";
                when x"145E" => data <= "00000";
                when x"145F" => data <= "11010";
                when x"1460" => data <= "00000";
                when x"1461" => data <= "00110";
                when x"1462" => data <= "00110";
                when x"1463" => data <= "00000";
                when x"1464" => data <= "00110";
                when x"1465" => data <= "00110";
                when x"1466" => data <= "11111";
                when x"1467" => data <= "00110";
                when x"1468" => data <= "01111";
                when x"1469" => data <= "10011";
                when x"146A" => data <= "00000";
                when x"146B" => data <= "00000";
                when x"146C" => data <= "00000";
                when x"146D" => data <= "00110";
                when x"146E" => data <= "00000";
                when x"146F" => data <= "00110";
                when x"1470" => data <= "01000";
                when x"1471" => data <= "00000";
                when x"1472" => data <= "00000";
                when x"1473" => data <= "00000";
                when x"1474" => data <= "00000";
                when x"1475" => data <= "00000";
                when x"1476" => data <= "01011";
                when x"1477" => data <= "00110";
                when x"1478" => data <= "00000";
                when x"1479" => data <= "00110";
                when x"147A" => data <= "00110";
                when x"147B" => data <= "00000";
                when x"147C" => data <= "00000";
                when x"147D" => data <= "00110";
                when x"147E" => data <= "00000";
                when x"147F" => data <= "00110";
                when x"1480" => data <= "00110";
                when x"1481" => data <= "00000";
                when x"1482" => data <= "00110";
                when x"1483" => data <= "00000";
                when x"1484" => data <= "00000";
                when x"1485" => data <= "00000";
                when x"1486" => data <= "00001";
                when x"1487" => data <= "00000";
                when x"1488" => data <= "00000";
                when x"1489" => data <= "00110";
                when x"148A" => data <= "00110";
                when x"148B" => data <= "00110";
                when x"148C" => data <= "00000";
                when x"148D" => data <= "00110";
                when x"148E" => data <= "00110";
                when x"148F" => data <= "00000";
                when x"1490" => data <= "00110";
                when x"1491" => data <= "00000";
                when x"1492" => data <= "11111";
                when x"1493" => data <= "00000";
                when x"1494" => data <= "00000";
                when x"1495" => data <= "00000";
                when x"1496" => data <= "00110";
                when x"1497" => data <= "00000";
                when x"1498" => data <= "00110";
                when x"1499" => data <= "00100";
                when x"149A" => data <= "00110";
                when x"149B" => data <= "10111";
                when x"149C" => data <= "00110";
                when x"149D" => data <= "00110";
                when x"149E" => data <= "00110";
                when x"149F" => data <= "00110";
                when x"14A0" => data <= "00000";
                when x"14A1" => data <= "00000";
                when x"14A2" => data <= "00110";
                when x"14A3" => data <= "00110";
                when x"14A4" => data <= "00000";
                when x"14A5" => data <= "00110";
                when x"14A6" => data <= "00000";
                when x"14A7" => data <= "00000";
                when x"14A8" => data <= "00000";
                when x"14A9" => data <= "00110";
                when x"14AA" => data <= "00000";
                when x"14AB" => data <= "00000";
                when x"14AC" => data <= "00110";
                when x"14AD" => data <= "00110";
                when x"14AE" => data <= "10111";
                when x"14AF" => data <= "00011";
                when x"14B0" => data <= "10101";
                when x"14B1" => data <= "00110";
                when x"14B2" => data <= "00000";
                when x"14B3" => data <= "01001";
                when x"14B4" => data <= "00110";
                when x"14B5" => data <= "00110";
                when x"14B6" => data <= "10111";
                when x"14B7" => data <= "00110";
                when x"14B8" => data <= "00110";
                when x"14B9" => data <= "00000";
                when x"14BA" => data <= "11101";
                when x"14BB" => data <= "01010";
                when x"14BC" => data <= "00110";
                when x"14BD" => data <= "00000";
                when x"14BE" => data <= "11000";
                when x"14BF" => data <= "00110";
                when x"14C0" => data <= "00110";
                when x"14C1" => data <= "00110";
                when x"14C2" => data <= "00000";
                when x"14C3" => data <= "00000";
                when x"14C4" => data <= "00110";
                when x"14C5" => data <= "00111";
                when x"14C6" => data <= "00000";
                when x"14C7" => data <= "00110";
                when x"14C8" => data <= "00000";
                when x"14C9" => data <= "00000";
                when x"14CA" => data <= "00110";
                when x"14CB" => data <= "00101";
                when x"14CC" => data <= "00110";
                when x"14CD" => data <= "00110";
                when x"14CE" => data <= "00000";
                when x"14CF" => data <= "00000";
                when x"14D0" => data <= "00000";
                when x"14D1" => data <= "00110";
                when x"14D2" => data <= "01001";
                when x"14D3" => data <= "00000";
                when x"14D4" => data <= "00110";
                when x"14D5" => data <= "00110";
                when x"14D6" => data <= "00110";
                when x"14D7" => data <= "11111";
                when x"14D8" => data <= "00000";
                when x"14D9" => data <= "00110";
                when x"14DA" => data <= "00110";
                when x"14DB" => data <= "00000";
                when x"14DC" => data <= "00000";
                when x"14DD" => data <= "00110";
                when x"14DE" => data <= "00110";
                when x"14DF" => data <= "00000";
                when x"14E0" => data <= "00110";
                when x"14E1" => data <= "00110";
                when x"14E2" => data <= "00110";
                when x"14E3" => data <= "00000";
                when x"14E4" => data <= "00000";
                when x"14E5" => data <= "00000";
                when x"14E6" => data <= "00110";
                when x"14E7" => data <= "11100";
                when x"14E8" => data <= "11001";
                when x"14E9" => data <= "00110";
                when x"14EA" => data <= "00110";
                when x"14EB" => data <= "11101";
                when x"14EC" => data <= "00000";
                when x"14ED" => data <= "00000";
                when x"14EE" => data <= "11111";
                when x"14EF" => data <= "00000";
                when x"14F0" => data <= "00110";
                when x"14F1" => data <= "00000";
                when x"14F2" => data <= "00110";
                when x"14F3" => data <= "00000";
                when x"14F4" => data <= "11111";
                when x"14F5" => data <= "00110";
                when x"14F6" => data <= "01010";
                when x"14F7" => data <= "00000";
                when x"14F8" => data <= "00110";
                when x"14F9" => data <= "00001";
                when x"14FA" => data <= "00110";
                when x"14FB" => data <= "10111";
                when x"14FC" => data <= "00110";
                when x"14FD" => data <= "00000";
                when x"14FE" => data <= "00000";
                when x"14FF" => data <= "00000";
                when x"1500" => data <= "00110";
                when x"1501" => data <= "00110";
                when x"1502" => data <= "00110";
                when x"1503" => data <= "01011";
                when x"1504" => data <= "00000";
                when x"1505" => data <= "00000";
                when x"1506" => data <= "00000";
                when x"1507" => data <= "00110";
                when x"1508" => data <= "00000";
                when x"1509" => data <= "00000";
                when x"150A" => data <= "00110";
                when x"150B" => data <= "00000";
                when x"150C" => data <= "00110";
                when x"150D" => data <= "00110";
                when x"150E" => data <= "00000";
                when x"150F" => data <= "11010";
                when x"1510" => data <= "00110";
                when x"1511" => data <= "00110";
                when x"1512" => data <= "00110";
                when x"1513" => data <= "00000";
                when x"1514" => data <= "00110";
                when x"1515" => data <= "10011";
                when x"1516" => data <= "00110";
                when x"1517" => data <= "00000";
                when x"1518" => data <= "00000";
                when x"1519" => data <= "00000";
                when x"151A" => data <= "00110";
                when x"151B" => data <= "00000";
                when x"151C" => data <= "00000";
                when x"151D" => data <= "01111";
                when x"151E" => data <= "00000";
                when x"151F" => data <= "00110";
                when x"1520" => data <= "00100";
                when x"1521" => data <= "00110";
                when x"1522" => data <= "01101";
                when x"1523" => data <= "00000";
                when x"1524" => data <= "11001";
                when x"1525" => data <= "00110";
                when x"1526" => data <= "00110";
                when x"1527" => data <= "00000";
                when x"1528" => data <= "00000";
                when x"1529" => data <= "01001";
                when x"152A" => data <= "00110";
                when x"152B" => data <= "00000";
                when x"152C" => data <= "00000";
                when x"152D" => data <= "00000";
                when x"152E" => data <= "01011";
                when x"152F" => data <= "00000";
                when x"1530" => data <= "10011";
                when x"1531" => data <= "00000";
                when x"1532" => data <= "00000";
                when x"1533" => data <= "00000";
                when x"1534" => data <= "00000";
                when x"1535" => data <= "00000";
                when x"1536" => data <= "00110";
                when x"1537" => data <= "00110";
                when x"1538" => data <= "00110";
                when x"1539" => data <= "00000";
                when x"153A" => data <= "00110";
                when x"153B" => data <= "00000";
                when x"153C" => data <= "00110";
                when x"153D" => data <= "00000";
                when x"153E" => data <= "00110";
                when x"153F" => data <= "00110";
                when x"1540" => data <= "10011";
                when x"1541" => data <= "00110";
                when x"1542" => data <= "00000";
                when x"1543" => data <= "00000";
                when x"1544" => data <= "00110";
                when x"1545" => data <= "00110";
                when x"1546" => data <= "00000";
                when x"1547" => data <= "00110";
                when x"1548" => data <= "00110";
                when x"1549" => data <= "00110";
                when x"154A" => data <= "01011";
                when x"154B" => data <= "00010";
                when x"154C" => data <= "00110";
                when x"154D" => data <= "00000";
                when x"154E" => data <= "10110";
                when x"154F" => data <= "00110";
                when x"1550" => data <= "10010";
                when x"1551" => data <= "00110";
                when x"1552" => data <= "00000";
                when x"1553" => data <= "00110";
                when x"1554" => data <= "00000";
                when x"1555" => data <= "00000";
                when x"1556" => data <= "00000";
                when x"1557" => data <= "00000";
                when x"1558" => data <= "10001";
                when x"1559" => data <= "01101";
                when x"155A" => data <= "00110";
                when x"155B" => data <= "11001";
                when x"155C" => data <= "01011";
                when x"155D" => data <= "00011";
                when x"155E" => data <= "00000";
                when x"155F" => data <= "00000";
                when x"1560" => data <= "00110";
                when x"1561" => data <= "01111";
                when x"1562" => data <= "00000";
                when x"1563" => data <= "00000";
                when x"1564" => data <= "00000";
                when x"1565" => data <= "00000";
                when x"1566" => data <= "00000";
                when x"1567" => data <= "00110";
                when x"1568" => data <= "01011";
                when x"1569" => data <= "01100";
                when x"156A" => data <= "00000";
                when x"156B" => data <= "11011";
                when x"156C" => data <= "00000";
                when x"156D" => data <= "01101";
                when x"156E" => data <= "00110";
                when x"156F" => data <= "00000";
                when x"1570" => data <= "00000";
                when x"1571" => data <= "00000";
                when x"1572" => data <= "01001";
                when x"1573" => data <= "01000";
                when x"1574" => data <= "11001";
                when x"1575" => data <= "01011";
                when x"1576" => data <= "00110";
                when x"1577" => data <= "00110";
                when x"1578" => data <= "00000";
                when x"1579" => data <= "00000";
                when x"157A" => data <= "00000";
                when x"157B" => data <= "11000";
                when x"157C" => data <= "00110";
                when x"157D" => data <= "00000";
                when x"157E" => data <= "00000";
                when x"157F" => data <= "00000";
                when x"1580" => data <= "00110";
                when x"1581" => data <= "00000";
                when x"1582" => data <= "00000";
                when x"1583" => data <= "11110";
                when x"1584" => data <= "00000";
                when x"1585" => data <= "00110";
                when x"1586" => data <= "00000";
                when x"1587" => data <= "00000";
                when x"1588" => data <= "00110";
                when x"1589" => data <= "00000";
                when x"158A" => data <= "00000";
                when x"158B" => data <= "11111";
                when x"158C" => data <= "00110";
                when x"158D" => data <= "10111";
                when x"158E" => data <= "00110";
                when x"158F" => data <= "00000";
                when x"1590" => data <= "00000";
                when x"1591" => data <= "00110";
                when x"1592" => data <= "00110";
                when x"1593" => data <= "11100";
                when x"1594" => data <= "00000";
                when x"1595" => data <= "00000";
                when x"1596" => data <= "00110";
                when x"1597" => data <= "00110";
                when x"1598" => data <= "00000";
                when x"1599" => data <= "00000";
                when x"159A" => data <= "00000";
                when x"159B" => data <= "00110";
                when x"159C" => data <= "00000";
                when x"159D" => data <= "00110";
                when x"159E" => data <= "00000";
                when x"159F" => data <= "00000";
                when x"15A0" => data <= "00110";
                when x"15A1" => data <= "00110";
                when x"15A2" => data <= "00011";
                when x"15A3" => data <= "11011";
                when x"15A4" => data <= "00000";
                when x"15A5" => data <= "00000";
                when x"15A6" => data <= "00000";
                when x"15A7" => data <= "00110";
                when x"15A8" => data <= "00000";
                when x"15A9" => data <= "00110";
                when x"15AA" => data <= "00110";
                when x"15AB" => data <= "00000";
                when x"15AC" => data <= "00000";
                when x"15AD" => data <= "00110";
                when x"15AE" => data <= "00110";
                when x"15AF" => data <= "00000";
                when x"15B0" => data <= "00110";
                when x"15B1" => data <= "10000";
                when x"15B2" => data <= "00000";
                when x"15B3" => data <= "00000";
                when x"15B4" => data <= "00000";
                when x"15B5" => data <= "01001";
                when x"15B6" => data <= "00000";
                when x"15B7" => data <= "00110";
                when x"15B8" => data <= "00000";
                when x"15B9" => data <= "00010";
                when x"15BA" => data <= "00110";
                when x"15BB" => data <= "00000";
                when x"15BC" => data <= "00000";
                when x"15BD" => data <= "00110";
                when x"15BE" => data <= "00000";
                when x"15BF" => data <= "00000";
                when x"15C0" => data <= "00000";
                when x"15C1" => data <= "00110";
                when x"15C2" => data <= "00000";
                when x"15C3" => data <= "00000";
                when x"15C4" => data <= "00110";
                when x"15C5" => data <= "10100";
                when x"15C6" => data <= "00000";
                when x"15C7" => data <= "11110";
                when x"15C8" => data <= "00110";
                when x"15C9" => data <= "01111";
                when x"15CA" => data <= "00110";
                when x"15CB" => data <= "00110";
                when x"15CC" => data <= "00110";
                when x"15CD" => data <= "00000";
                when x"15CE" => data <= "00000";
                when x"15CF" => data <= "00000";
                when x"15D0" => data <= "00110";
                when x"15D1" => data <= "00000";
                when x"15D2" => data <= "00000";
                when x"15D3" => data <= "01110";
                when x"15D4" => data <= "00000";
                when x"15D5" => data <= "00110";
                when x"15D6" => data <= "00000";
                when x"15D7" => data <= "00000";
                when x"15D8" => data <= "00000";
                when x"15D9" => data <= "00110";
                when x"15DA" => data <= "00000";
                when x"15DB" => data <= "00000";
                when x"15DC" => data <= "00000";
                when x"15DD" => data <= "00000";
                when x"15DE" => data <= "00110";
                when x"15DF" => data <= "00110";
                when x"15E0" => data <= "00000";
                when x"15E1" => data <= "01011";
                when x"15E2" => data <= "10010";
                when x"15E3" => data <= "00110";
                when x"15E4" => data <= "00101";
                when x"15E5" => data <= "00000";
                when x"15E6" => data <= "00110";
                when x"15E7" => data <= "00000";
                when x"15E8" => data <= "00110";
                when x"15E9" => data <= "00110";
                when x"15EA" => data <= "00000";
                when x"15EB" => data <= "11110";
                when x"15EC" => data <= "01010";
                when x"15ED" => data <= "00000";
                when x"15EE" => data <= "00110";
                when x"15EF" => data <= "00110";
                when x"15F0" => data <= "00000";
                when x"15F1" => data <= "01111";
                when x"15F2" => data <= "00110";
                when x"15F3" => data <= "00000";
                when x"15F4" => data <= "00110";
                when x"15F5" => data <= "00000";
                when x"15F6" => data <= "01011";
                when x"15F7" => data <= "10011";
                when x"15F8" => data <= "11100";
                when x"15F9" => data <= "00000";
                when x"15FA" => data <= "00110";
                when x"15FB" => data <= "00000";
                when x"15FC" => data <= "00110";
                when x"15FD" => data <= "00110";
                when x"15FE" => data <= "00110";
                when x"15FF" => data <= "00110";
                when x"1600" => data <= "00110";
                when x"1601" => data <= "00110";
                when x"1602" => data <= "00000";
                when x"1603" => data <= "00000";
                when x"1604" => data <= "11011";
                when x"1605" => data <= "00000";
                when x"1606" => data <= "00000";
                when x"1607" => data <= "00000";
                when x"1608" => data <= "00110";
                when x"1609" => data <= "00000";
                when x"160A" => data <= "00000";
                when x"160B" => data <= "00000";
                when x"160C" => data <= "00000";
                when x"160D" => data <= "10111";
                when x"160E" => data <= "00000";
                when x"160F" => data <= "10011";
                when x"1610" => data <= "00000";
                when x"1611" => data <= "00000";
                when x"1612" => data <= "00110";
                when x"1613" => data <= "00000";
                when x"1614" => data <= "00110";
                when x"1615" => data <= "00000";
                when x"1616" => data <= "00000";
                when x"1617" => data <= "00000";
                when x"1618" => data <= "10011";
                when x"1619" => data <= "00110";
                when x"161A" => data <= "00000";
                when x"161B" => data <= "00110";
                when x"161C" => data <= "00110";
                when x"161D" => data <= "00110";
                when x"161E" => data <= "00000";
                when x"161F" => data <= "11000";
                when x"1620" => data <= "01101";
                when x"1621" => data <= "00000";
                when x"1622" => data <= "00000";
                when x"1623" => data <= "00110";
                when x"1624" => data <= "00000";
                when x"1625" => data <= "00000";
                when x"1626" => data <= "00000";
                when x"1627" => data <= "00000";
                when x"1628" => data <= "00110";
                when x"1629" => data <= "00011";
                when x"162A" => data <= "00000";
                when x"162B" => data <= "00110";
                when x"162C" => data <= "00000";
                when x"162D" => data <= "00000";
                when x"162E" => data <= "11101";
                when x"162F" => data <= "01011";
                when x"1630" => data <= "00110";
                when x"1631" => data <= "00110";
                when x"1632" => data <= "00000";
                when x"1633" => data <= "00110";
                when x"1634" => data <= "00110";
                when x"1635" => data <= "00110";
                when x"1636" => data <= "01011";
                when x"1637" => data <= "00000";
                when x"1638" => data <= "00000";
                when x"1639" => data <= "00110";
                when x"163A" => data <= "00000";
                when x"163B" => data <= "00110";
                when x"163C" => data <= "00000";
                when x"163D" => data <= "00110";
                when x"163E" => data <= "11100";
                when x"163F" => data <= "00000";
                when x"1640" => data <= "01111";
                when x"1641" => data <= "00000";
                when x"1642" => data <= "00000";
                when x"1643" => data <= "00110";
                when x"1644" => data <= "00110";
                when x"1645" => data <= "00000";
                when x"1646" => data <= "00110";
                when x"1647" => data <= "00000";
                when x"1648" => data <= "00000";
                when x"1649" => data <= "00000";
                when x"164A" => data <= "00110";
                when x"164B" => data <= "00000";
                when x"164C" => data <= "00000";
                when x"164D" => data <= "01011";
                when x"164E" => data <= "00000";
                when x"164F" => data <= "01100";
                when x"1650" => data <= "00110";
                when x"1651" => data <= "00110";
                when x"1652" => data <= "00001";
                when x"1653" => data <= "00000";
                when x"1654" => data <= "00000";
                when x"1655" => data <= "00000";
                when x"1656" => data <= "00000";
                when x"1657" => data <= "00101";
                when x"1658" => data <= "00110";
                when x"1659" => data <= "00110";
                when x"165A" => data <= "00000";
                when x"165B" => data <= "01101";
                when x"165C" => data <= "00110";
                when x"165D" => data <= "00000";
                when x"165E" => data <= "01111";
                when x"165F" => data <= "00000";
                when x"1660" => data <= "00000";
                when x"1661" => data <= "00000";
                when x"1662" => data <= "00110";
                when x"1663" => data <= "00000";
                when x"1664" => data <= "00110";
                when x"1665" => data <= "00110";
                when x"1666" => data <= "00000";
                when x"1667" => data <= "00000";
                when x"1668" => data <= "01100";
                when x"1669" => data <= "11111";
                when x"166A" => data <= "00000";
                when x"166B" => data <= "00000";
                when x"166C" => data <= "00110";
                when x"166D" => data <= "00011";
                when x"166E" => data <= "00110";
                when x"166F" => data <= "10101";
                when x"1670" => data <= "00110";
                when x"1671" => data <= "11111";
                when x"1672" => data <= "00000";
                when x"1673" => data <= "01111";
                when x"1674" => data <= "00000";
                when x"1675" => data <= "10001";
                when x"1676" => data <= "00110";
                when x"1677" => data <= "00000";
                when x"1678" => data <= "00110";
                when x"1679" => data <= "01100";
                when x"167A" => data <= "00110";
                when x"167B" => data <= "10001";
                when x"167C" => data <= "00000";
                when x"167D" => data <= "00110";
                when x"167E" => data <= "00000";
                when x"167F" => data <= "00110";
                when x"1680" => data <= "00000";
                when x"1681" => data <= "00101";
                when x"1682" => data <= "00000";
                when x"1683" => data <= "00000";
                when x"1684" => data <= "11110";
                when x"1685" => data <= "00110";
                when x"1686" => data <= "00000";
                when x"1687" => data <= "11001";
                when x"1688" => data <= "01101";
                when x"1689" => data <= "11001";
                when x"168A" => data <= "00000";
                when x"168B" => data <= "00000";
                when x"168C" => data <= "00110";
                when x"168D" => data <= "00000";
                when x"168E" => data <= "00110";
                when x"168F" => data <= "00000";
                when x"1690" => data <= "00110";
                when x"1691" => data <= "00110";
                when x"1692" => data <= "00110";
                when x"1693" => data <= "00110";
                when x"1694" => data <= "00000";
                when x"1695" => data <= "00000";
                when x"1696" => data <= "11111";
                when x"1697" => data <= "00110";
                when x"1698" => data <= "00000";
                when x"1699" => data <= "00110";
                when x"169A" => data <= "01101";
                when x"169B" => data <= "00000";
                when x"169C" => data <= "00000";
                when x"169D" => data <= "00000";
                when x"169E" => data <= "10011";
                when x"169F" => data <= "00110";
                when x"16A0" => data <= "00000";
                when x"16A1" => data <= "10011";
                when x"16A2" => data <= "00101";
                when x"16A3" => data <= "00010";
                when x"16A4" => data <= "00000";
                when x"16A5" => data <= "00110";
                when x"16A6" => data <= "00000";
                when x"16A7" => data <= "00000";
                when x"16A8" => data <= "11001";
                when x"16A9" => data <= "01001";
                when x"16AA" => data <= "11000";
                when x"16AB" => data <= "00110";
                when x"16AC" => data <= "00110";
                when x"16AD" => data <= "00110";
                when x"16AE" => data <= "01101";
                when x"16AF" => data <= "01101";
                when x"16B0" => data <= "00000";
                when x"16B1" => data <= "10000";
                when x"16B2" => data <= "11001";
                when x"16B3" => data <= "00000";
                when x"16B4" => data <= "00000";
                when x"16B5" => data <= "00000";
                when x"16B6" => data <= "00110";
                when x"16B7" => data <= "00110";
                when x"16B8" => data <= "00110";
                when x"16B9" => data <= "00110";
                when x"16BA" => data <= "00000";
                when x"16BB" => data <= "00110";
                when x"16BC" => data <= "00000";
                when x"16BD" => data <= "00000";
                when x"16BE" => data <= "00000";
                when x"16BF" => data <= "00110";
                when x"16C0" => data <= "00110";
                when x"16C1" => data <= "00110";
                when x"16C2" => data <= "00000";
                when x"16C3" => data <= "00000";
                when x"16C4" => data <= "00000";
                when x"16C5" => data <= "00110";
                when x"16C6" => data <= "00000";
                when x"16C7" => data <= "00110";
                when x"16C8" => data <= "01111";
                when x"16C9" => data <= "00000";
                when x"16CA" => data <= "00000";
                when x"16CB" => data <= "00110";
                when x"16CC" => data <= "00000";
                when x"16CD" => data <= "00000";
                when x"16CE" => data <= "00011";
                when x"16CF" => data <= "00000";
                when x"16D0" => data <= "00110";
                when x"16D1" => data <= "00100";
                when x"16D2" => data <= "00110";
                when x"16D3" => data <= "00110";
                when x"16D4" => data <= "01011";
                when x"16D5" => data <= "00000";
                when x"16D6" => data <= "00110";
                when x"16D7" => data <= "00000";
                when x"16D8" => data <= "00110";
                when x"16D9" => data <= "11001";
                when x"16DA" => data <= "10001";
                when x"16DB" => data <= "00000";
                when x"16DC" => data <= "00110";
                when x"16DD" => data <= "00000";
                when x"16DE" => data <= "00000";
                when x"16DF" => data <= "00000";
                when x"16E0" => data <= "00110";
                when x"16E1" => data <= "00000";
                when x"16E2" => data <= "00110";
                when x"16E3" => data <= "00000";
                when x"16E4" => data <= "01011";
                when x"16E5" => data <= "11101";
                when x"16E6" => data <= "00110";
                when x"16E7" => data <= "00110";
                when x"16E8" => data <= "00110";
                when x"16E9" => data <= "00110";
                when x"16EA" => data <= "11111";
                when x"16EB" => data <= "00110";
                when x"16EC" => data <= "00000";
                when x"16ED" => data <= "00000";
                when x"16EE" => data <= "00110";
                when x"16EF" => data <= "00110";
                when x"16F0" => data <= "00110";
                when x"16F1" => data <= "00000";
                when x"16F2" => data <= "00110";
                when x"16F3" => data <= "00000";
                when x"16F4" => data <= "00110";
                when x"16F5" => data <= "00000";
                when x"16F6" => data <= "00000";
                when x"16F7" => data <= "00110";
                when x"16F8" => data <= "00110";
                when x"16F9" => data <= "00110";
                when x"16FA" => data <= "00000";
                when x"16FB" => data <= "00110";
                when x"16FC" => data <= "00000";
                when x"16FD" => data <= "10001";
                when x"16FE" => data <= "00000";
                when x"16FF" => data <= "00110";
                when x"1700" => data <= "00000";
                when x"1701" => data <= "00000";
                when x"1702" => data <= "00110";
                when x"1703" => data <= "00000";
                when x"1704" => data <= "00000";
                when x"1705" => data <= "00000";
                when x"1706" => data <= "00110";
                when x"1707" => data <= "00000";
                when x"1708" => data <= "00000";
                when x"1709" => data <= "00000";
                when x"170A" => data <= "00110";
                when x"170B" => data <= "01011";
                when x"170C" => data <= "00000";
                when x"170D" => data <= "00110";
                when x"170E" => data <= "10111";
                when x"170F" => data <= "00110";
                when x"1710" => data <= "00000";
                when x"1711" => data <= "00110";
                when x"1712" => data <= "00110";
                when x"1713" => data <= "00110";
                when x"1714" => data <= "00110";
                when x"1715" => data <= "10101";
                when x"1716" => data <= "10010";
                when x"1717" => data <= "00000";
                when x"1718" => data <= "00110";
                when x"1719" => data <= "00000";
                when x"171A" => data <= "00110";
                when x"171B" => data <= "00000";
                when x"171C" => data <= "00000";
                when x"171D" => data <= "00000";
                when x"171E" => data <= "00000";
                when x"171F" => data <= "10011";
                when x"1720" => data <= "00000";
                when x"1721" => data <= "00110";
                when x"1722" => data <= "11100";
                when x"1723" => data <= "00110";
                when x"1724" => data <= "11011";
                when x"1725" => data <= "00110";
                when x"1726" => data <= "00000";
                when x"1727" => data <= "00000";
                when x"1728" => data <= "00110";
                when x"1729" => data <= "11100";
                when x"172A" => data <= "00110";
                when x"172B" => data <= "00110";
                when x"172C" => data <= "00110";
                when x"172D" => data <= "11001";
                when x"172E" => data <= "00010";
                when x"172F" => data <= "01011";
                when x"1730" => data <= "00000";
                when x"1731" => data <= "00110";
                when x"1732" => data <= "00110";
                when x"1733" => data <= "00000";
                when x"1734" => data <= "00000";
                when x"1735" => data <= "00000";
                when x"1736" => data <= "00110";
                when x"1737" => data <= "00110";
                when x"1738" => data <= "00000";
                when x"1739" => data <= "00110";
                when x"173A" => data <= "00000";
                when x"173B" => data <= "00000";
                when x"173C" => data <= "00000";
                when x"173D" => data <= "00000";
                when x"173E" => data <= "00110";
                when x"173F" => data <= "00000";
                when x"1740" => data <= "00000";
                when x"1741" => data <= "00110";
                when x"1742" => data <= "00110";
                when x"1743" => data <= "00000";
                when x"1744" => data <= "00110";
                when x"1745" => data <= "00000";
                when x"1746" => data <= "00110";
                when x"1747" => data <= "00110";
                when x"1748" => data <= "00101";
                when x"1749" => data <= "11010";
                when x"174A" => data <= "00000";
                when x"174B" => data <= "11101";
                when x"174C" => data <= "10011";
                when x"174D" => data <= "10100";
                when x"174E" => data <= "10011";
                when x"174F" => data <= "00110";
                when x"1750" => data <= "00000";
                when x"1751" => data <= "00000";
                when x"1752" => data <= "00000";
                when x"1753" => data <= "00110";
                when x"1754" => data <= "00000";
                when x"1755" => data <= "01011";
                when x"1756" => data <= "00110";
                when x"1757" => data <= "00110";
                when x"1758" => data <= "00110";
                when x"1759" => data <= "00000";
                when x"175A" => data <= "00000";
                when x"175B" => data <= "00110";
                when x"175C" => data <= "00000";
                when x"175D" => data <= "00110";
                when x"175E" => data <= "00000";
                when x"175F" => data <= "01101";
                when x"1760" => data <= "10011";
                when x"1761" => data <= "00110";
                when x"1762" => data <= "00110";
                when x"1763" => data <= "00110";
                when x"1764" => data <= "01011";
                when x"1765" => data <= "01110";
                when x"1766" => data <= "00000";
                when x"1767" => data <= "00000";
                when x"1768" => data <= "00110";
                when x"1769" => data <= "00000";
                when x"176A" => data <= "00000";
                when x"176B" => data <= "00000";
                when x"176C" => data <= "10110";
                when x"176D" => data <= "00110";
                when x"176E" => data <= "00110";
                when x"176F" => data <= "00110";
                when x"1770" => data <= "00000";
                when x"1771" => data <= "00000";
                when x"1772" => data <= "00011";
                when x"1773" => data <= "00110";
                when x"1774" => data <= "00000";
                when x"1775" => data <= "00011";
                when x"1776" => data <= "00001";
                when x"1777" => data <= "00000";
                when x"1778" => data <= "00000";
                when x"1779" => data <= "00000";
                when x"177A" => data <= "00000";
                when x"177B" => data <= "00110";
                when x"177C" => data <= "00000";
                when x"177D" => data <= "00110";
                when x"177E" => data <= "00110";
                when x"177F" => data <= "11011";
                when x"1780" => data <= "00110";
                when x"1781" => data <= "01101";
                when x"1782" => data <= "00110";
                when x"1783" => data <= "00110";
                when x"1784" => data <= "00110";
                when x"1785" => data <= "10011";
                when x"1786" => data <= "00110";
                when x"1787" => data <= "00000";
                when x"1788" => data <= "00000";
                when x"1789" => data <= "00110";
                when x"178A" => data <= "10000";
                when x"178B" => data <= "00000";
                when x"178C" => data <= "00000";
                when x"178D" => data <= "00110";
                when x"178E" => data <= "00000";
                when x"178F" => data <= "00111";
                when x"1790" => data <= "00000";
                when x"1791" => data <= "00000";
                when x"1792" => data <= "00110";
                when x"1793" => data <= "00110";
                when x"1794" => data <= "00000";
                when x"1795" => data <= "10000";
                when x"1796" => data <= "00000";
                when x"1797" => data <= "00110";
                when x"1798" => data <= "00000";
                when x"1799" => data <= "00000";
                when x"179A" => data <= "10100";
                when x"179B" => data <= "00110";
                when x"179C" => data <= "01011";
                when x"179D" => data <= "11001";
                when x"179E" => data <= "00110";
                when x"179F" => data <= "00110";
                when x"17A0" => data <= "01011";
                when x"17A1" => data <= "00011";
                when x"17A2" => data <= "00000";
                when x"17A3" => data <= "00000";
                when x"17A4" => data <= "00110";
                when x"17A5" => data <= "00110";
                when x"17A6" => data <= "01011";
                when x"17A7" => data <= "10010";
                when x"17A8" => data <= "00000";
                when x"17A9" => data <= "00110";
                when x"17AA" => data <= "00000";
                when x"17AB" => data <= "00110";
                when x"17AC" => data <= "00110";
                when x"17AD" => data <= "11001";
                when x"17AE" => data <= "00000";
                when x"17AF" => data <= "10011";
                when x"17B0" => data <= "00000";
                when x"17B1" => data <= "00110";
                when x"17B2" => data <= "00000";
                when x"17B3" => data <= "00000";
                when x"17B4" => data <= "00000";
                when x"17B5" => data <= "00110";
                when x"17B6" => data <= "00000";
                when x"17B7" => data <= "11100";
                when x"17B8" => data <= "00110";
                when x"17B9" => data <= "00110";
                when x"17BA" => data <= "00000";
                when x"17BB" => data <= "00000";
                when x"17BC" => data <= "00110";
                when x"17BD" => data <= "00100";
                when x"17BE" => data <= "00000";
                when x"17BF" => data <= "00000";
                when x"17C0" => data <= "00110";
                when x"17C1" => data <= "00000";
                when x"17C2" => data <= "00110";
                when x"17C3" => data <= "00110";
                when x"17C4" => data <= "00110";
                when x"17C5" => data <= "00000";
                when x"17C6" => data <= "10101";
                when x"17C7" => data <= "00110";
                when x"17C8" => data <= "00000";
                when x"17C9" => data <= "00110";
                when x"17CA" => data <= "00000";
                when x"17CB" => data <= "01110";
                when x"17CC" => data <= "11001";
                when x"17CD" => data <= "00110";
                when x"17CE" => data <= "00110";
                when x"17CF" => data <= "00110";
                when x"17D0" => data <= "11001";
                when x"17D1" => data <= "00000";
                when x"17D2" => data <= "00110";
                when x"17D3" => data <= "11101";
                when x"17D4" => data <= "10011";
                when x"17D5" => data <= "00110";
                when x"17D6" => data <= "01011";
                when x"17D7" => data <= "00110";
                when x"17D8" => data <= "00110";
                when x"17D9" => data <= "00110";
                when x"17DA" => data <= "00000";
                when x"17DB" => data <= "00100";
                when x"17DC" => data <= "10011";
                when x"17DD" => data <= "10010";
                when x"17DE" => data <= "00000";
                when x"17DF" => data <= "00000";
                when x"17E0" => data <= "10100";
                when x"17E1" => data <= "00110";
                when x"17E2" => data <= "00110";
                when x"17E3" => data <= "00000";
                when x"17E4" => data <= "00000";
                when x"17E5" => data <= "01011";
                when x"17E6" => data <= "00110";
                when x"17E7" => data <= "00000";
                when x"17E8" => data <= "00000";
                when x"17E9" => data <= "00110";
                when x"17EA" => data <= "00000";
                when x"17EB" => data <= "00000";
                when x"17EC" => data <= "11100";
                when x"17ED" => data <= "00110";
                when x"17EE" => data <= "00000";
                when x"17EF" => data <= "11010";
                when x"17F0" => data <= "00000";
                when x"17F1" => data <= "00000";
                when x"17F2" => data <= "10001";
                when x"17F3" => data <= "00000";
                when x"17F4" => data <= "00000";
                when x"17F5" => data <= "00110";
                when x"17F6" => data <= "00110";
                when x"17F7" => data <= "00110";
                when x"17F8" => data <= "00000";
                when x"17F9" => data <= "00000";
                when x"17FA" => data <= "00000";
                when x"17FB" => data <= "00000";
                when x"17FC" => data <= "00000";
                when x"17FD" => data <= "00110";
                when x"17FE" => data <= "00110";
                when x"17FF" => data <= "00110";
                when x"1800" => data <= "00000";
                when x"1801" => data <= "00000";
                when x"1802" => data <= "00110";
                when x"1803" => data <= "00110";
                when x"1804" => data <= "00000";
                when x"1805" => data <= "00110";
                when x"1806" => data <= "01111";
                when x"1807" => data <= "00000";
                when x"1808" => data <= "00000";
                when x"1809" => data <= "01110";
                when x"180A" => data <= "11001";
                when x"180B" => data <= "00110";
                when x"180C" => data <= "00110";
                when x"180D" => data <= "00000";
                when x"180E" => data <= "11001";
                when x"180F" => data <= "00110";
                when x"1810" => data <= "00000";
                when x"1811" => data <= "01100";
                when x"1812" => data <= "11001";
                when x"1813" => data <= "00110";
                when x"1814" => data <= "01101";
                when x"1815" => data <= "00110";
                when x"1816" => data <= "01101";
                when x"1817" => data <= "01011";
                when x"1818" => data <= "00000";
                when x"1819" => data <= "00110";
                when x"181A" => data <= "00000";
                when x"181B" => data <= "00011";
                when x"181C" => data <= "00000";
                when x"181D" => data <= "00000";
                when x"181E" => data <= "00110";
                when x"181F" => data <= "00000";
                when x"1820" => data <= "00000";
                when x"1821" => data <= "00110";
                when x"1822" => data <= "00000";
                when x"1823" => data <= "11110";
                when x"1824" => data <= "00110";
                when x"1825" => data <= "00000";
                when x"1826" => data <= "00000";
                when x"1827" => data <= "00110";
                when x"1828" => data <= "00000";
                when x"1829" => data <= "01100";
                when x"182A" => data <= "10011";
                when x"182B" => data <= "00110";
                when x"182C" => data <= "00110";
                when x"182D" => data <= "00110";
                when x"182E" => data <= "00110";
                when x"182F" => data <= "00110";
                when x"1830" => data <= "00000";
                when x"1831" => data <= "00110";
                when x"1832" => data <= "00000";
                when x"1833" => data <= "00110";
                when x"1834" => data <= "00110";
                when x"1835" => data <= "00000";
                when x"1836" => data <= "00000";
                when x"1837" => data <= "00110";
                when x"1838" => data <= "00110";
                when x"1839" => data <= "11000";
                when x"183A" => data <= "00110";
                when x"183B" => data <= "00110";
                when x"183C" => data <= "00000";
                when x"183D" => data <= "00110";
                when x"183E" => data <= "00000";
                when x"183F" => data <= "00000";
                when x"1840" => data <= "00000";
                when x"1841" => data <= "10101";
                when x"1842" => data <= "00000";
                when x"1843" => data <= "00110";
                when x"1844" => data <= "00110";
                when x"1845" => data <= "00110";
                when x"1846" => data <= "00000";
                when x"1847" => data <= "00000";
                when x"1848" => data <= "00000";
                when x"1849" => data <= "00000";
                when x"184A" => data <= "00000";
                when x"184B" => data <= "00110";
                when x"184C" => data <= "01101";
                when x"184D" => data <= "00000";
                when x"184E" => data <= "00110";
                when x"184F" => data <= "00000";
                when x"1850" => data <= "00110";
                when x"1851" => data <= "00000";
                when x"1852" => data <= "00000";
                when x"1853" => data <= "00110";
                when x"1854" => data <= "00110";
                when x"1855" => data <= "00110";
                when x"1856" => data <= "10011";
                when x"1857" => data <= "01010";
                when x"1858" => data <= "00110";
                when x"1859" => data <= "00110";
                when x"185A" => data <= "00000";
                when x"185B" => data <= "01011";
                when x"185C" => data <= "01010";
                when x"185D" => data <= "00000";
                when x"185E" => data <= "00000";
                when x"185F" => data <= "00000";
                when x"1860" => data <= "00110";
                when x"1861" => data <= "00110";
                when x"1862" => data <= "00000";
                when x"1863" => data <= "00110";
                when x"1864" => data <= "11010";
                when x"1865" => data <= "00110";
                when x"1866" => data <= "01101";
                when x"1867" => data <= "00110";
                when x"1868" => data <= "00110";
                when x"1869" => data <= "00000";
                when x"186A" => data <= "00000";
                when x"186B" => data <= "00000";
                when x"186C" => data <= "00000";
                when x"186D" => data <= "00000";
                when x"186E" => data <= "00110";
                when x"186F" => data <= "00000";
                when x"1870" => data <= "00000";
                when x"1871" => data <= "00110";
                when x"1872" => data <= "00110";
                when x"1873" => data <= "00110";
                when x"1874" => data <= "00110";
                when x"1875" => data <= "00000";
                when x"1876" => data <= "00110";
                when x"1877" => data <= "00000";
                when x"1878" => data <= "01100";
                when x"1879" => data <= "00000";
                when x"187A" => data <= "00010";
                when x"187B" => data <= "00110";
                when x"187C" => data <= "00110";
                when x"187D" => data <= "00000";
                when x"187E" => data <= "00110";
                when x"187F" => data <= "01110";
                when x"1880" => data <= "00110";
                when x"1881" => data <= "00000";
                when x"1882" => data <= "00000";
                when x"1883" => data <= "00001";
                when x"1884" => data <= "00000";
                when x"1885" => data <= "00110";
                when x"1886" => data <= "00010";
                when x"1887" => data <= "00110";
                when x"1888" => data <= "00000";
                when x"1889" => data <= "00110";
                when x"188A" => data <= "00011";
                when x"188B" => data <= "00110";
                when x"188C" => data <= "10000";
                when x"188D" => data <= "00110";
                when x"188E" => data <= "00000";
                when x"188F" => data <= "00110";
                when x"1890" => data <= "00110";
                when x"1891" => data <= "00000";
                when x"1892" => data <= "00110";
                when x"1893" => data <= "00000";
                when x"1894" => data <= "11011";
                when x"1895" => data <= "00000";
                when x"1896" => data <= "00000";
                when x"1897" => data <= "01011";
                when x"1898" => data <= "00000";
                when x"1899" => data <= "00110";
                when x"189A" => data <= "00110";
                when x"189B" => data <= "10110";
                when x"189C" => data <= "00110";
                when x"189D" => data <= "00000";
                when x"189E" => data <= "00000";
                when x"189F" => data <= "11111";
                when x"18A0" => data <= "00110";
                when x"18A1" => data <= "00100";
                when x"18A2" => data <= "00000";
                when x"18A3" => data <= "01101";
                when x"18A4" => data <= "00000";
                when x"18A5" => data <= "10001";
                when x"18A6" => data <= "00000";
                when x"18A7" => data <= "00110";
                when x"18A8" => data <= "11111";
                when x"18A9" => data <= "00110";
                when x"18AA" => data <= "00110";
                when x"18AB" => data <= "10111";
                when x"18AC" => data <= "00000";
                when x"18AD" => data <= "00110";
                when x"18AE" => data <= "00110";
                when x"18AF" => data <= "00110";
                when x"18B0" => data <= "10100";
                when x"18B1" => data <= "00000";
                when x"18B2" => data <= "00000";
                when x"18B3" => data <= "00110";
                when x"18B4" => data <= "10000";
                when x"18B5" => data <= "10010";
                when x"18B6" => data <= "00000";
                when x"18B7" => data <= "00000";
                when x"18B8" => data <= "00001";
                when x"18B9" => data <= "00110";
                when x"18BA" => data <= "00000";
                when x"18BB" => data <= "10100";
                when x"18BC" => data <= "00110";
                when x"18BD" => data <= "00110";
                when x"18BE" => data <= "00110";
                when x"18BF" => data <= "00000";
                when x"18C0" => data <= "00110";
                when x"18C1" => data <= "00001";
                when x"18C2" => data <= "00000";
                when x"18C3" => data <= "00110";
                when x"18C4" => data <= "00110";
                when x"18C5" => data <= "10000";
                when x"18C6" => data <= "00000";
                when x"18C7" => data <= "00000";
                when x"18C8" => data <= "00000";
                when x"18C9" => data <= "01010";
                when x"18CA" => data <= "00000";
                when x"18CB" => data <= "10000";
                when x"18CC" => data <= "11001";
                when x"18CD" => data <= "00000";
                when x"18CE" => data <= "11001";
                when x"18CF" => data <= "00000";
                when x"18D0" => data <= "00110";
                when x"18D1" => data <= "00110";
                when x"18D2" => data <= "00001";
                when x"18D3" => data <= "00000";
                when x"18D4" => data <= "00000";
                when x"18D5" => data <= "00000";
                when x"18D6" => data <= "00000";
                when x"18D7" => data <= "00110";
                when x"18D8" => data <= "00110";
                when x"18D9" => data <= "00000";
                when x"18DA" => data <= "00010";
                when x"18DB" => data <= "00000";
                when x"18DC" => data <= "00110";
                when x"18DD" => data <= "00000";
                when x"18DE" => data <= "10100";
                when x"18DF" => data <= "00000";
                when x"18E0" => data <= "00000";
                when x"18E1" => data <= "00110";
                when x"18E2" => data <= "00000";
                when x"18E3" => data <= "00110";
                when x"18E4" => data <= "00110";
                when x"18E5" => data <= "00110";
                when x"18E6" => data <= "00000";
                when x"18E7" => data <= "00110";
                when x"18E8" => data <= "00110";
                when x"18E9" => data <= "00110";
                when x"18EA" => data <= "00000";
                when x"18EB" => data <= "11101";
                when x"18EC" => data <= "10101";
                when x"18ED" => data <= "00000";
                when x"18EE" => data <= "00110";
                when x"18EF" => data <= "00110";
                when x"18F0" => data <= "00000";
                when x"18F1" => data <= "00000";
                when x"18F2" => data <= "01110";
                when x"18F3" => data <= "11001";
                when x"18F4" => data <= "00000";
                when x"18F5" => data <= "00001";
                when x"18F6" => data <= "00000";
                when x"18F7" => data <= "00000";
                when x"18F8" => data <= "00000";
                when x"18F9" => data <= "00000";
                when x"18FA" => data <= "00000";
                when x"18FB" => data <= "00110";
                when x"18FC" => data <= "00110";
                when x"18FD" => data <= "00110";
                when x"18FE" => data <= "00000";
                when x"18FF" => data <= "00000";
                when x"1900" => data <= "01000";
                when x"1901" => data <= "00000";
                when x"1902" => data <= "00000";
                when x"1903" => data <= "10110";
                when x"1904" => data <= "00000";
                when x"1905" => data <= "00110";
                when x"1906" => data <= "00000";
                when x"1907" => data <= "00110";
                when x"1908" => data <= "00110";
                when x"1909" => data <= "00110";
                when x"190A" => data <= "00000";
                when x"190B" => data <= "00110";
                when x"190C" => data <= "01111";
                when x"190D" => data <= "00110";
                when x"190E" => data <= "00110";
                when x"190F" => data <= "00110";
                when x"1910" => data <= "00000";
                when x"1911" => data <= "00110";
                when x"1912" => data <= "00000";
                when x"1913" => data <= "00110";
                when x"1914" => data <= "00110";
                when x"1915" => data <= "00110";
                when x"1916" => data <= "00000";
                when x"1917" => data <= "00110";
                when x"1918" => data <= "00000";
                when x"1919" => data <= "00110";
                when x"191A" => data <= "00000";
                when x"191B" => data <= "00110";
                when x"191C" => data <= "00110";
                when x"191D" => data <= "00110";
                when x"191E" => data <= "10011";
                when x"191F" => data <= "00110";
                when x"1920" => data <= "11111";
                when x"1921" => data <= "00110";
                when x"1922" => data <= "00000";
                when x"1923" => data <= "00000";
                when x"1924" => data <= "00110";
                when x"1925" => data <= "00110";
                when x"1926" => data <= "00010";
                when x"1927" => data <= "00000";
                when x"1928" => data <= "00110";
                when x"1929" => data <= "00110";
                when x"192A" => data <= "01111";
                when x"192B" => data <= "00000";
                when x"192C" => data <= "00000";
                when x"192D" => data <= "11111";
                when x"192E" => data <= "00000";
                when x"192F" => data <= "00110";
                when x"1930" => data <= "00110";
                when x"1931" => data <= "00000";
                when x"1932" => data <= "10011";
                when x"1933" => data <= "00000";
                when x"1934" => data <= "00101";
                when x"1935" => data <= "11100";
                when x"1936" => data <= "00110";
                when x"1937" => data <= "00110";
                when x"1938" => data <= "00000";
                when x"1939" => data <= "01100";
                when x"193A" => data <= "00110";
                when x"193B" => data <= "00110";
                when x"193C" => data <= "01101";
                when x"193D" => data <= "00000";
                when x"193E" => data <= "01110";
                when x"193F" => data <= "10010";
                when x"1940" => data <= "00000";
                when x"1941" => data <= "00110";
                when x"1942" => data <= "00000";
                when x"1943" => data <= "00110";
                when x"1944" => data <= "00000";
                when x"1945" => data <= "10001";
                when x"1946" => data <= "00000";
                when x"1947" => data <= "00110";
                when x"1948" => data <= "00010";
                when x"1949" => data <= "00000";
                when x"194A" => data <= "11111";
                when x"194B" => data <= "00110";
                when x"194C" => data <= "00110";
                when x"194D" => data <= "00110";
                when x"194E" => data <= "00110";
                when x"194F" => data <= "00110";
                when x"1950" => data <= "00110";
                when x"1951" => data <= "00000";
                when x"1952" => data <= "00000";
                when x"1953" => data <= "00000";
                when x"1954" => data <= "10001";
                when x"1955" => data <= "00111";
                when x"1956" => data <= "00000";
                when x"1957" => data <= "00110";
                when x"1958" => data <= "00000";
                when x"1959" => data <= "00000";
                when x"195A" => data <= "00000";
                when x"195B" => data <= "00000";
                when x"195C" => data <= "00000";
                when x"195D" => data <= "00000";
                when x"195E" => data <= "00000";
                when x"195F" => data <= "00000";
                when x"1960" => data <= "00000";
                when x"1961" => data <= "00000";
                when x"1962" => data <= "00110";
                when x"1963" => data <= "10000";
                when x"1964" => data <= "10001";
                when x"1965" => data <= "00110";
                when x"1966" => data <= "00110";
                when x"1967" => data <= "00110";
                when x"1968" => data <= "00000";
                when x"1969" => data <= "01001";
                when x"196A" => data <= "00110";
                when x"196B" => data <= "00110";
                when x"196C" => data <= "00110";
                when x"196D" => data <= "00000";
                when x"196E" => data <= "10111";
                when x"196F" => data <= "00000";
                when x"1970" => data <= "00110";
                when x"1971" => data <= "00000";
                when x"1972" => data <= "00000";
                when x"1973" => data <= "11001";
                when x"1974" => data <= "00110";
                when x"1975" => data <= "11001";
                when x"1976" => data <= "01001";
                when x"1977" => data <= "00000";
                when x"1978" => data <= "00110";
                when x"1979" => data <= "00000";
                when x"197A" => data <= "00000";
                when x"197B" => data <= "01001";
                when x"197C" => data <= "01001";
                when x"197D" => data <= "00110";
                when x"197E" => data <= "11010";
                when x"197F" => data <= "10111";
                when x"1980" => data <= "00000";
                when x"1981" => data <= "01100";
                when x"1982" => data <= "00110";
                when x"1983" => data <= "00000";
                when x"1984" => data <= "01000";
                when x"1985" => data <= "00000";
                when x"1986" => data <= "00110";
                when x"1987" => data <= "00110";
                when x"1988" => data <= "00000";
                when x"1989" => data <= "00000";
                when x"198A" => data <= "00000";
                when x"198B" => data <= "00000";
                when x"198C" => data <= "00000";
                when x"198D" => data <= "00000";
                when x"198E" => data <= "00000";
                when x"198F" => data <= "00110";
                when x"1990" => data <= "00110";
                when x"1991" => data <= "00000";
                when x"1992" => data <= "00110";
                when x"1993" => data <= "00000";
                when x"1994" => data <= "00110";
                when x"1995" => data <= "00110";
                when x"1996" => data <= "00000";
                when x"1997" => data <= "00110";
                when x"1998" => data <= "00000";
                when x"1999" => data <= "10010";
                when x"199A" => data <= "00000";
                when x"199B" => data <= "01101";
                when x"199C" => data <= "00000";
                when x"199D" => data <= "00000";
                when x"199E" => data <= "11110";
                when x"199F" => data <= "00000";
                when x"19A0" => data <= "00000";
                when x"19A1" => data <= "01101";
                when x"19A2" => data <= "00000";
                when x"19A3" => data <= "01111";
                when x"19A4" => data <= "00110";
                when x"19A5" => data <= "00110";
                when x"19A6" => data <= "00110";
                when x"19A7" => data <= "11010";
                when x"19A8" => data <= "00000";
                when x"19A9" => data <= "00000";
                when x"19AA" => data <= "00110";
                when x"19AB" => data <= "11011";
                when x"19AC" => data <= "00110";
                when x"19AD" => data <= "00110";
                when x"19AE" => data <= "00000";
                when x"19AF" => data <= "00000";
                when x"19B0" => data <= "00000";
                when x"19B1" => data <= "00110";
                when x"19B2" => data <= "00110";
                when x"19B3" => data <= "00000";
                when x"19B4" => data <= "00000";
                when x"19B5" => data <= "00000";
                when x"19B6" => data <= "00000";
                when x"19B7" => data <= "00110";
                when x"19B8" => data <= "11100";
                when x"19B9" => data <= "00110";
                when x"19BA" => data <= "00000";
                when x"19BB" => data <= "00110";
                when x"19BC" => data <= "10111";
                when x"19BD" => data <= "00000";
                when x"19BE" => data <= "00000";
                when x"19BF" => data <= "00000";
                when x"19C0" => data <= "00110";
                when x"19C1" => data <= "00110";
                when x"19C2" => data <= "00000";
                when x"19C3" => data <= "00110";
                when x"19C4" => data <= "00110";
                when x"19C5" => data <= "00110";
                when x"19C6" => data <= "01011";
                when x"19C7" => data <= "11111";
                when x"19C8" => data <= "00110";
                when x"19C9" => data <= "00000";
                when x"19CA" => data <= "01101";
                when x"19CB" => data <= "00000";
                when x"19CC" => data <= "00000";
                when x"19CD" => data <= "00001";
                when x"19CE" => data <= "00000";
                when x"19CF" => data <= "00000";
                when x"19D0" => data <= "00000";
                when x"19D1" => data <= "00000";
                when x"19D2" => data <= "00000";
                when x"19D3" => data <= "01011";
                when x"19D4" => data <= "11100";
                when x"19D5" => data <= "00000";
                when x"19D6" => data <= "01011";
                when x"19D7" => data <= "00110";
                when x"19D8" => data <= "00000";
                when x"19D9" => data <= "00110";
                when x"19DA" => data <= "00110";
                when x"19DB" => data <= "00000";
                when x"19DC" => data <= "00000";
                when x"19DD" => data <= "00110";
                when x"19DE" => data <= "00110";
                when x"19DF" => data <= "00111";
                when x"19E0" => data <= "00000";
                when x"19E1" => data <= "00000";
                when x"19E2" => data <= "00010";
                when x"19E3" => data <= "00110";
                when x"19E4" => data <= "00000";
                when x"19E5" => data <= "00000";
                when x"19E6" => data <= "00110";
                when x"19E7" => data <= "00110";
                when x"19E8" => data <= "00110";
                when x"19E9" => data <= "00110";
                when x"19EA" => data <= "00000";
                when x"19EB" => data <= "00000";
                when x"19EC" => data <= "00110";
                when x"19ED" => data <= "00110";
                when x"19EE" => data <= "00000";
                when x"19EF" => data <= "11111";
                when x"19F0" => data <= "00110";
                when x"19F1" => data <= "00000";
                when x"19F2" => data <= "00000";
                when x"19F3" => data <= "00000";
                when x"19F4" => data <= "00110";
                when x"19F5" => data <= "00110";
                when x"19F6" => data <= "00110";
                when x"19F7" => data <= "00110";
                when x"19F8" => data <= "00000";
                when x"19F9" => data <= "00000";
                when x"19FA" => data <= "00000";
                when x"19FB" => data <= "00000";
                when x"19FC" => data <= "00001";
                when x"19FD" => data <= "01001";
                when x"19FE" => data <= "00000";
                when x"19FF" => data <= "00110";
                when x"1A00" => data <= "00110";
                when x"1A01" => data <= "00000";
                when x"1A02" => data <= "00000";
                when x"1A03" => data <= "00110";
                when x"1A04" => data <= "00000";
                when x"1A05" => data <= "00000";
                when x"1A06" => data <= "01010";
                when x"1A07" => data <= "00110";
                when x"1A08" => data <= "00110";
                when x"1A09" => data <= "00000";
                when x"1A0A" => data <= "00110";
                when x"1A0B" => data <= "00110";
                when x"1A0C" => data <= "00000";
                when x"1A0D" => data <= "00110";
                when x"1A0E" => data <= "00000";
                when x"1A0F" => data <= "00000";
                when x"1A10" => data <= "00110";
                when x"1A11" => data <= "10000";
                when x"1A12" => data <= "00110";
                when x"1A13" => data <= "00000";
                when x"1A14" => data <= "00110";
                when x"1A15" => data <= "00000";
                when x"1A16" => data <= "00110";
                when x"1A17" => data <= "00000";
                when x"1A18" => data <= "00000";
                when x"1A19" => data <= "00000";
                when x"1A1A" => data <= "00110";
                when x"1A1B" => data <= "11011";
                when x"1A1C" => data <= "00000";
                when x"1A1D" => data <= "01111";
                when x"1A1E" => data <= "00000";
                when x"1A1F" => data <= "00110";
                when x"1A20" => data <= "00110";
                when x"1A21" => data <= "00110";
                when x"1A22" => data <= "00110";
                when x"1A23" => data <= "10011";
                when x"1A24" => data <= "00111";
                when x"1A25" => data <= "00000";
                when x"1A26" => data <= "00000";
                when x"1A27" => data <= "00000";
                when x"1A28" => data <= "00000";
                when x"1A29" => data <= "00110";
                when x"1A2A" => data <= "01101";
                when x"1A2B" => data <= "00000";
                when x"1A2C" => data <= "00110";
                when x"1A2D" => data <= "00110";
                when x"1A2E" => data <= "00000";
                when x"1A2F" => data <= "00000";
                when x"1A30" => data <= "00000";
                when x"1A31" => data <= "00000";
                when x"1A32" => data <= "00000";
                when x"1A33" => data <= "00000";
                when x"1A34" => data <= "00000";
                when x"1A35" => data <= "00000";
                when x"1A36" => data <= "00000";
                when x"1A37" => data <= "00000";
                when x"1A38" => data <= "00110";
                when x"1A39" => data <= "10000";
                when x"1A3A" => data <= "00110";
                when x"1A3B" => data <= "00110";
                when x"1A3C" => data <= "11000";
                when x"1A3D" => data <= "00110";
                when x"1A3E" => data <= "00110";
                when x"1A3F" => data <= "10101";
                when x"1A40" => data <= "00000";
                when x"1A41" => data <= "00110";
                when x"1A42" => data <= "00110";
                when x"1A43" => data <= "01101";
                when x"1A44" => data <= "00000";
                when x"1A45" => data <= "00110";
                when x"1A46" => data <= "00000";
                when x"1A47" => data <= "00000";
                when x"1A48" => data <= "00000";
                when x"1A49" => data <= "01011";
                when x"1A4A" => data <= "00000";
                when x"1A4B" => data <= "00110";
                when x"1A4C" => data <= "01101";
                when x"1A4D" => data <= "00110";
                when x"1A4E" => data <= "00100";
                when x"1A4F" => data <= "00110";
                when x"1A50" => data <= "00101";
                when x"1A51" => data <= "00110";
                when x"1A52" => data <= "00000";
                when x"1A53" => data <= "00110";
                when x"1A54" => data <= "00000";
                when x"1A55" => data <= "01111";
                when x"1A56" => data <= "00000";
                when x"1A57" => data <= "01000";
                when x"1A58" => data <= "00000";
                when x"1A59" => data <= "00000";
                when x"1A5A" => data <= "00000";
                when x"1A5B" => data <= "00110";
                when x"1A5C" => data <= "00000";
                when x"1A5D" => data <= "10010";
                when x"1A5E" => data <= "00110";
                when x"1A5F" => data <= "01100";
                when x"1A60" => data <= "00100";
                when x"1A61" => data <= "00000";
                when x"1A62" => data <= "00110";
                when x"1A63" => data <= "00000";
                when x"1A64" => data <= "00110";
                when x"1A65" => data <= "00000";
                when x"1A66" => data <= "00110";
                when x"1A67" => data <= "00110";
                when x"1A68" => data <= "00000";
                when x"1A69" => data <= "00000";
                when x"1A6A" => data <= "00000";
                when x"1A6B" => data <= "00000";
                when x"1A6C" => data <= "00110";
                when x"1A6D" => data <= "00110";
                when x"1A6E" => data <= "00110";
                when x"1A6F" => data <= "00110";
                when x"1A70" => data <= "00000";
                when x"1A71" => data <= "01011";
                when x"1A72" => data <= "00110";
                when x"1A73" => data <= "00110";
                when x"1A74" => data <= "00110";
                when x"1A75" => data <= "00000";
                when x"1A76" => data <= "00000";
                when x"1A77" => data <= "01100";
                when x"1A78" => data <= "00110";
                when x"1A79" => data <= "10111";
                when x"1A7A" => data <= "00110";
                when x"1A7B" => data <= "01001";
                when x"1A7C" => data <= "00000";
                when x"1A7D" => data <= "11111";
                when x"1A7E" => data <= "00000";
                when x"1A7F" => data <= "00110";
                when x"1A80" => data <= "00110";
                when x"1A81" => data <= "00000";
                when x"1A82" => data <= "00000";
                when x"1A83" => data <= "00000";
                when x"1A84" => data <= "00000";
                when x"1A85" => data <= "01110";
                when x"1A86" => data <= "01011";
                when x"1A87" => data <= "00000";
                when x"1A88" => data <= "01010";
                when x"1A89" => data <= "00000";
                when x"1A8A" => data <= "00000";
                when x"1A8B" => data <= "00000";
                when x"1A8C" => data <= "11111";
                when x"1A8D" => data <= "00000";
                when x"1A8E" => data <= "00110";
                when x"1A8F" => data <= "00110";
                when x"1A90" => data <= "00110";
                when x"1A91" => data <= "00110";
                when x"1A92" => data <= "00110";
                when x"1A93" => data <= "00110";
                when x"1A94" => data <= "00000";
                when x"1A95" => data <= "00000";
                when x"1A96" => data <= "00000";
                when x"1A97" => data <= "00000";
                when x"1A98" => data <= "00110";
                when x"1A99" => data <= "00000";
                when x"1A9A" => data <= "11001";
                when x"1A9B" => data <= "00110";
                when x"1A9C" => data <= "00000";
                when x"1A9D" => data <= "10011";
                when x"1A9E" => data <= "00110";
                when x"1A9F" => data <= "00110";
                when x"1AA0" => data <= "00110";
                when x"1AA1" => data <= "00000";
                when x"1AA2" => data <= "00000";
                when x"1AA3" => data <= "00110";
                when x"1AA4" => data <= "00000";
                when x"1AA5" => data <= "00000";
                when x"1AA6" => data <= "01011";
                when x"1AA7" => data <= "00000";
                when x"1AA8" => data <= "00110";
                when x"1AA9" => data <= "00000";
                when x"1AAA" => data <= "00000";
                when x"1AAB" => data <= "00000";
                when x"1AAC" => data <= "00110";
                when x"1AAD" => data <= "00110";
                when x"1AAE" => data <= "00110";
                when x"1AAF" => data <= "11111";
                when x"1AB0" => data <= "00110";
                when x"1AB1" => data <= "00011";
                when x"1AB2" => data <= "00000";
                when x"1AB3" => data <= "11110";
                when x"1AB4" => data <= "01011";
                when x"1AB5" => data <= "00110";
                when x"1AB6" => data <= "00000";
                when x"1AB7" => data <= "01111";
                when x"1AB8" => data <= "00000";
                when x"1AB9" => data <= "11100";
                when x"1ABA" => data <= "00000";
                when x"1ABB" => data <= "10000";
                when x"1ABC" => data <= "00000";
                when x"1ABD" => data <= "00000";
                when x"1ABE" => data <= "00000";
                when x"1ABF" => data <= "00110";
                when x"1AC0" => data <= "00000";
                when x"1AC1" => data <= "00000";
                when x"1AC2" => data <= "00110";
                when x"1AC3" => data <= "10101";
                when x"1AC4" => data <= "00110";
                when x"1AC5" => data <= "00000";
                when x"1AC6" => data <= "00110";
                when x"1AC7" => data <= "00000";
                when x"1AC8" => data <= "00110";
                when x"1AC9" => data <= "00000";
                when x"1ACA" => data <= "11011";
                when x"1ACB" => data <= "00000";
                when x"1ACC" => data <= "00110";
                when x"1ACD" => data <= "00110";
                when x"1ACE" => data <= "00000";
                when x"1ACF" => data <= "00000";
                when x"1AD0" => data <= "00000";
                when x"1AD1" => data <= "10100";
                when x"1AD2" => data <= "00110";
                when x"1AD3" => data <= "00000";
                when x"1AD4" => data <= "00000";
                when x"1AD5" => data <= "00000";
                when x"1AD6" => data <= "00000";
                when x"1AD7" => data <= "00000";
                when x"1AD8" => data <= "10001";
                when x"1AD9" => data <= "01011";
                when x"1ADA" => data <= "00110";
                when x"1ADB" => data <= "11001";
                when x"1ADC" => data <= "00110";
                when x"1ADD" => data <= "00110";
                when x"1ADE" => data <= "00110";
                when x"1ADF" => data <= "00000";
                when x"1AE0" => data <= "00000";
                when x"1AE1" => data <= "00000";
                when x"1AE2" => data <= "00000";
                when x"1AE3" => data <= "00000";
                when x"1AE4" => data <= "00110";
                when x"1AE5" => data <= "00000";
                when x"1AE6" => data <= "01111";
                when x"1AE7" => data <= "00110";
                when x"1AE8" => data <= "00000";
                when x"1AE9" => data <= "01101";
                when x"1AEA" => data <= "00000";
                when x"1AEB" => data <= "00110";
                when x"1AEC" => data <= "00000";
                when x"1AED" => data <= "00110";
                when x"1AEE" => data <= "00000";
                when x"1AEF" => data <= "00000";
                when x"1AF0" => data <= "00000";
                when x"1AF1" => data <= "00000";
                when x"1AF2" => data <= "00110";
                when x"1AF3" => data <= "00110";
                when x"1AF4" => data <= "00110";
                when x"1AF5" => data <= "00000";
                when x"1AF6" => data <= "00000";
                when x"1AF7" => data <= "00110";
                when x"1AF8" => data <= "01010";
                when x"1AF9" => data <= "00000";
                when x"1AFA" => data <= "00110";
                when x"1AFB" => data <= "00000";
                when x"1AFC" => data <= "00110";
                when x"1AFD" => data <= "00000";
                when x"1AFE" => data <= "00110";
                when x"1AFF" => data <= "01001";
                when x"1B00" => data <= "11111";
                when x"1B01" => data <= "00000";
                when x"1B02" => data <= "11000";
                when x"1B03" => data <= "01101";
                when x"1B04" => data <= "00110";
                when x"1B05" => data <= "00000";
                when x"1B06" => data <= "11001";
                when x"1B07" => data <= "00110";
                when x"1B08" => data <= "00000";
                when x"1B09" => data <= "00110";
                when x"1B0A" => data <= "00000";
                when x"1B0B" => data <= "11010";
                when x"1B0C" => data <= "00000";
                when x"1B0D" => data <= "00000";
                when x"1B0E" => data <= "00000";
                when x"1B0F" => data <= "00000";
                when x"1B10" => data <= "00000";
                when x"1B11" => data <= "00000";
                when x"1B12" => data <= "11111";
                when x"1B13" => data <= "11111";
                when x"1B14" => data <= "00110";
                when x"1B15" => data <= "00000";
                when x"1B16" => data <= "01001";
                when x"1B17" => data <= "00110";
                when x"1B18" => data <= "00110";
                when x"1B19" => data <= "00000";
                when x"1B1A" => data <= "00110";
                when x"1B1B" => data <= "00000";
                when x"1B1C" => data <= "00110";
                when x"1B1D" => data <= "00000";
                when x"1B1E" => data <= "00000";
                when x"1B1F" => data <= "00000";
                when x"1B20" => data <= "11001";
                when x"1B21" => data <= "00110";
                when x"1B22" => data <= "10001";
                when x"1B23" => data <= "00000";
                when x"1B24" => data <= "00110";
                when x"1B25" => data <= "00000";
                when x"1B26" => data <= "00000";
                when x"1B27" => data <= "00110";
                when x"1B28" => data <= "00000";
                when x"1B29" => data <= "10001";
                when x"1B2A" => data <= "00110";
                when x"1B2B" => data <= "00110";
                when x"1B2C" => data <= "01011";
                when x"1B2D" => data <= "00000";
                when x"1B2E" => data <= "00000";
                when x"1B2F" => data <= "00000";
                when x"1B30" => data <= "10000";
                when x"1B31" => data <= "00000";
                when x"1B32" => data <= "00000";
                when x"1B33" => data <= "00110";
                when x"1B34" => data <= "00110";
                when x"1B35" => data <= "10111";
                when x"1B36" => data <= "00110";
                when x"1B37" => data <= "00000";
                when x"1B38" => data <= "00110";
                when x"1B39" => data <= "00000";
                when x"1B3A" => data <= "10001";
                when x"1B3B" => data <= "00000";
                when x"1B3C" => data <= "00000";
                when x"1B3D" => data <= "10000";
                when x"1B3E" => data <= "00000";
                when x"1B3F" => data <= "01000";
                when x"1B40" => data <= "00000";
                when x"1B41" => data <= "00110";
                when x"1B42" => data <= "00000";
                when x"1B43" => data <= "00000";
                when x"1B44" => data <= "00000";
                when x"1B45" => data <= "00000";
                when x"1B46" => data <= "00000";
                when x"1B47" => data <= "00110";
                when x"1B48" => data <= "00000";
                when x"1B49" => data <= "00110";
                when x"1B4A" => data <= "00000";
                when x"1B4B" => data <= "00110";
                when x"1B4C" => data <= "00110";
                when x"1B4D" => data <= "00000";
                when x"1B4E" => data <= "00000";
                when x"1B4F" => data <= "00110";
                when x"1B50" => data <= "01010";
                when x"1B51" => data <= "00110";
                when x"1B52" => data <= "00110";
                when x"1B53" => data <= "00110";
                when x"1B54" => data <= "10010";
                when x"1B55" => data <= "00000";
                when x"1B56" => data <= "00110";
                when x"1B57" => data <= "00110";
                when x"1B58" => data <= "00110";
                when x"1B59" => data <= "00110";
                when x"1B5A" => data <= "00000";
                when x"1B5B" => data <= "00000";
                when x"1B5C" => data <= "00110";
                when x"1B5D" => data <= "00110";
                when x"1B5E" => data <= "00000";
                when x"1B5F" => data <= "00110";
                when x"1B60" => data <= "01010";
                when x"1B61" => data <= "00110";
                when x"1B62" => data <= "00000";
                when x"1B63" => data <= "00110";
                when x"1B64" => data <= "00000";
                when x"1B65" => data <= "00110";
                when x"1B66" => data <= "00110";
                when x"1B67" => data <= "00000";
                when x"1B68" => data <= "00000";
                when x"1B69" => data <= "00000";
                when x"1B6A" => data <= "10100";
                when x"1B6B" => data <= "00000";
                when x"1B6C" => data <= "00110";
                when x"1B6D" => data <= "00110";
                when x"1B6E" => data <= "00000";
                when x"1B6F" => data <= "00000";
                when x"1B70" => data <= "10100";
                when x"1B71" => data <= "00000";
                when x"1B72" => data <= "00000";
                when x"1B73" => data <= "11010";
                when x"1B74" => data <= "01101";
                when x"1B75" => data <= "11111";
                when x"1B76" => data <= "00000";
                when x"1B77" => data <= "01101";
                when x"1B78" => data <= "01001";
                when x"1B79" => data <= "00110";
                when x"1B7A" => data <= "00110";
                when x"1B7B" => data <= "00000";
                when x"1B7C" => data <= "00000";
                when x"1B7D" => data <= "00110";
                when x"1B7E" => data <= "00000";
                when x"1B7F" => data <= "00000";
                when x"1B80" => data <= "01101";
                when x"1B81" => data <= "00000";
                when x"1B82" => data <= "00000";
                when x"1B83" => data <= "00000";
                when x"1B84" => data <= "00000";
                when x"1B85" => data <= "10010";
                when x"1B86" => data <= "00000";
                when x"1B87" => data <= "00000";
                when x"1B88" => data <= "00000";
                when x"1B89" => data <= "00000";
                when x"1B8A" => data <= "00110";
                when x"1B8B" => data <= "11011";
                when x"1B8C" => data <= "00110";
                when x"1B8D" => data <= "10110";
                when x"1B8E" => data <= "00110";
                when x"1B8F" => data <= "00110";
                when x"1B90" => data <= "00110";
                when x"1B91" => data <= "00011";
                when x"1B92" => data <= "00000";
                when x"1B93" => data <= "00110";
                when x"1B94" => data <= "00000";
                when x"1B95" => data <= "00110";
                when x"1B96" => data <= "00110";
                when x"1B97" => data <= "00110";
                when x"1B98" => data <= "00000";
                when x"1B99" => data <= "00000";
                when x"1B9A" => data <= "00110";
                when x"1B9B" => data <= "00110";
                when x"1B9C" => data <= "00000";
                when x"1B9D" => data <= "00110";
                when x"1B9E" => data <= "00000";
                when x"1B9F" => data <= "00110";
                when x"1BA0" => data <= "00110";
                when x"1BA1" => data <= "10011";
                when x"1BA2" => data <= "01100";
                when x"1BA3" => data <= "00110";
                when x"1BA4" => data <= "00110";
                when x"1BA5" => data <= "11101";
                when x"1BA6" => data <= "00110";
                when x"1BA7" => data <= "00110";
                when x"1BA8" => data <= "00000";
                when x"1BA9" => data <= "00000";
                when x"1BAA" => data <= "00000";
                when x"1BAB" => data <= "00000";
                when x"1BAC" => data <= "00110";
                when x"1BAD" => data <= "00110";
                when x"1BAE" => data <= "10100";
                when x"1BAF" => data <= "00110";
                when x"1BB0" => data <= "00110";
                when x"1BB1" => data <= "00000";
                when x"1BB2" => data <= "00110";
                when x"1BB3" => data <= "00000";
                when x"1BB4" => data <= "00110";
                when x"1BB5" => data <= "00110";
                when x"1BB6" => data <= "11001";
                when x"1BB7" => data <= "00110";
                when x"1BB8" => data <= "01101";
                when x"1BB9" => data <= "00000";
                when x"1BBA" => data <= "00110";
                when x"1BBB" => data <= "00000";
                when x"1BBC" => data <= "01110";
                when x"1BBD" => data <= "00000";
                when x"1BBE" => data <= "01011";
                when x"1BBF" => data <= "00110";
                when x"1BC0" => data <= "00000";
                when x"1BC1" => data <= "00110";
                when x"1BC2" => data <= "00000";
                when x"1BC3" => data <= "11000";
                when x"1BC4" => data <= "00000";
                when x"1BC5" => data <= "01011";
                when x"1BC6" => data <= "00000";
                when x"1BC7" => data <= "00000";
                when x"1BC8" => data <= "10101";
                when x"1BC9" => data <= "00000";
                when x"1BCA" => data <= "00000";
                when x"1BCB" => data <= "00110";
                when x"1BCC" => data <= "00000";
                when x"1BCD" => data <= "00000";
                when x"1BCE" => data <= "00000";
                when x"1BCF" => data <= "00110";
                when x"1BD0" => data <= "01011";
                when x"1BD1" => data <= "11101";
                when x"1BD2" => data <= "00000";
                when x"1BD3" => data <= "00010";
                when x"1BD4" => data <= "00000";
                when x"1BD5" => data <= "00110";
                when x"1BD6" => data <= "00011";
                when x"1BD7" => data <= "00000";
                when x"1BD8" => data <= "00000";
                when x"1BD9" => data <= "00000";
                when x"1BDA" => data <= "00110";
                when x"1BDB" => data <= "00110";
                when x"1BDC" => data <= "00110";
                when x"1BDD" => data <= "00000";
                when x"1BDE" => data <= "00000";
                when x"1BDF" => data <= "10101";
                when x"1BE0" => data <= "00110";
                when x"1BE1" => data <= "00000";
                when x"1BE2" => data <= "00000";
                when x"1BE3" => data <= "00000";
                when x"1BE4" => data <= "00000";
                when x"1BE5" => data <= "00110";
                when x"1BE6" => data <= "00000";
                when x"1BE7" => data <= "00000";
                when x"1BE8" => data <= "00000";
                when x"1BE9" => data <= "00110";
                when x"1BEA" => data <= "01110";
                when x"1BEB" => data <= "00000";
                when x"1BEC" => data <= "01011";
                when x"1BED" => data <= "11110";
                when x"1BEE" => data <= "00000";
                when x"1BEF" => data <= "00000";
                when x"1BF0" => data <= "00001";
                when x"1BF1" => data <= "00110";
                when x"1BF2" => data <= "00000";
                when x"1BF3" => data <= "11001";
                when x"1BF4" => data <= "00110";
                when x"1BF5" => data <= "00000";
                when x"1BF6" => data <= "01110";
                when x"1BF7" => data <= "00000";
                when x"1BF8" => data <= "00110";
                when x"1BF9" => data <= "10100";
                when x"1BFA" => data <= "00000";
                when x"1BFB" => data <= "00110";
                when x"1BFC" => data <= "00000";
                when x"1BFD" => data <= "00000";
                when x"1BFE" => data <= "00110";
                when x"1BFF" => data <= "00110";
                when x"1C00" => data <= "00110";
                when x"1C01" => data <= "00001";
                when x"1C02" => data <= "00110";
                when x"1C03" => data <= "00000";
                when x"1C04" => data <= "00110";
                when x"1C05" => data <= "00000";
                when x"1C06" => data <= "00110";
                when x"1C07" => data <= "00110";
                when x"1C08" => data <= "11001";
                when x"1C09" => data <= "00001";
                when x"1C0A" => data <= "00000";
                when x"1C0B" => data <= "10001";
                when x"1C0C" => data <= "10101";
                when x"1C0D" => data <= "00000";
                when x"1C0E" => data <= "10111";
                when x"1C0F" => data <= "00110";
                when x"1C10" => data <= "00110";
                when x"1C11" => data <= "00000";
                when x"1C12" => data <= "10101";
                when x"1C13" => data <= "10101";
                when x"1C14" => data <= "00110";
                when x"1C15" => data <= "00000";
                when x"1C16" => data <= "00000";
                when x"1C17" => data <= "00110";
                when x"1C18" => data <= "00110";
                when x"1C19" => data <= "00000";
                when x"1C1A" => data <= "01010";
                when x"1C1B" => data <= "00000";
                when x"1C1C" => data <= "00110";
                when x"1C1D" => data <= "00000";
                when x"1C1E" => data <= "10111";
                when x"1C1F" => data <= "00110";
                when x"1C20" => data <= "01001";
                when x"1C21" => data <= "00110";
                when x"1C22" => data <= "00000";
                when x"1C23" => data <= "11110";
                when x"1C24" => data <= "00000";
                when x"1C25" => data <= "01101";
                when x"1C26" => data <= "00000";
                when x"1C27" => data <= "00110";
                when x"1C28" => data <= "00110";
                when x"1C29" => data <= "00110";
                when x"1C2A" => data <= "00000";
                when x"1C2B" => data <= "11101";
                when x"1C2C" => data <= "00000";
                when x"1C2D" => data <= "00000";
                when x"1C2E" => data <= "00000";
                when x"1C2F" => data <= "00000";
                when x"1C30" => data <= "00110";
                when x"1C31" => data <= "00110";
                when x"1C32" => data <= "00011";
                when x"1C33" => data <= "00000";
                when x"1C34" => data <= "00111";
                when x"1C35" => data <= "11011";
                when x"1C36" => data <= "00111";
                when x"1C37" => data <= "11101";
                when x"1C38" => data <= "00000";
                when x"1C39" => data <= "10000";
                when x"1C3A" => data <= "00000";
                when x"1C3B" => data <= "01101";
                when x"1C3C" => data <= "00000";
                when x"1C3D" => data <= "00110";
                when x"1C3E" => data <= "00000";
                when x"1C3F" => data <= "00000";
                when x"1C40" => data <= "00110";
                when x"1C41" => data <= "00000";
                when x"1C42" => data <= "01010";
                when x"1C43" => data <= "00110";
                when x"1C44" => data <= "00000";
                when x"1C45" => data <= "00110";
                when x"1C46" => data <= "00110";
                when x"1C47" => data <= "00110";
                when x"1C48" => data <= "00000";
                when x"1C49" => data <= "00110";
                when x"1C4A" => data <= "00110";
                when x"1C4B" => data <= "00110";
                when x"1C4C" => data <= "01011";
                when x"1C4D" => data <= "01100";
                when x"1C4E" => data <= "00000";
                when x"1C4F" => data <= "00110";
                when x"1C50" => data <= "00000";
                when x"1C51" => data <= "00000";
                when x"1C52" => data <= "10100";
                when x"1C53" => data <= "11001";
                when x"1C54" => data <= "00110";
                when x"1C55" => data <= "00110";
                when x"1C56" => data <= "00110";
                when x"1C57" => data <= "00110";
                when x"1C58" => data <= "00000";
                when x"1C59" => data <= "00000";
                when x"1C5A" => data <= "00110";
                when x"1C5B" => data <= "10001";
                when x"1C5C" => data <= "11110";
                when x"1C5D" => data <= "00110";
                when x"1C5E" => data <= "00000";
                when x"1C5F" => data <= "00110";
                when x"1C60" => data <= "01011";
                when x"1C61" => data <= "00110";
                when x"1C62" => data <= "00110";
                when x"1C63" => data <= "00110";
                when x"1C64" => data <= "00110";
                when x"1C65" => data <= "11100";
                when x"1C66" => data <= "00000";
                when x"1C67" => data <= "00110";
                when x"1C68" => data <= "10001";
                when x"1C69" => data <= "00000";
                when x"1C6A" => data <= "00110";
                when x"1C6B" => data <= "00000";
                when x"1C6C" => data <= "11010";
                when x"1C6D" => data <= "00000";
                when x"1C6E" => data <= "00110";
                when x"1C6F" => data <= "00110";
                when x"1C70" => data <= "00110";
                when x"1C71" => data <= "10101";
                when x"1C72" => data <= "00110";
                when x"1C73" => data <= "01110";
                when x"1C74" => data <= "00110";
                when x"1C75" => data <= "00000";
                when x"1C76" => data <= "00110";
                when x"1C77" => data <= "00110";
                when x"1C78" => data <= "00110";
                when x"1C79" => data <= "00110";
                when x"1C7A" => data <= "00111";
                when x"1C7B" => data <= "00000";
                when x"1C7C" => data <= "00000";
                when x"1C7D" => data <= "00110";
                when x"1C7E" => data <= "00110";
                when x"1C7F" => data <= "00110";
                when x"1C80" => data <= "00000";
                when x"1C81" => data <= "00000";
                when x"1C82" => data <= "00000";
                when x"1C83" => data <= "00000";
                when x"1C84" => data <= "00000";
                when x"1C85" => data <= "10011";
                when x"1C86" => data <= "00110";
                when x"1C87" => data <= "01011";
                when x"1C88" => data <= "00000";
                when x"1C89" => data <= "00110";
                when x"1C8A" => data <= "00110";
                when x"1C8B" => data <= "00000";
                when x"1C8C" => data <= "10001";
                when x"1C8D" => data <= "00000";
                when x"1C8E" => data <= "01011";
                when x"1C8F" => data <= "00000";
                when x"1C90" => data <= "11011";
                when x"1C91" => data <= "00110";
                when x"1C92" => data <= "01011";
                when x"1C93" => data <= "00000";
                when x"1C94" => data <= "01101";
                when x"1C95" => data <= "11110";
                when x"1C96" => data <= "00110";
                when x"1C97" => data <= "00110";
                when x"1C98" => data <= "00110";
                when x"1C99" => data <= "00000";
                when x"1C9A" => data <= "00000";
                when x"1C9B" => data <= "00110";
                when x"1C9C" => data <= "00001";
                when x"1C9D" => data <= "00110";
                when x"1C9E" => data <= "00110";
                when x"1C9F" => data <= "00000";
                when x"1CA0" => data <= "00110";
                when x"1CA1" => data <= "00110";
                when x"1CA2" => data <= "00000";
                when x"1CA3" => data <= "00110";
                when x"1CA4" => data <= "00110";
                when x"1CA5" => data <= "00000";
                when x"1CA6" => data <= "00000";
                when x"1CA7" => data <= "00000";
                when x"1CA8" => data <= "00011";
                when x"1CA9" => data <= "00110";
                when x"1CAA" => data <= "00000";
                when x"1CAB" => data <= "00110";
                when x"1CAC" => data <= "00110";
                when x"1CAD" => data <= "00110";
                when x"1CAE" => data <= "00000";
                when x"1CAF" => data <= "00000";
                when x"1CB0" => data <= "10100";
                when x"1CB1" => data <= "00000";
                when x"1CB2" => data <= "00000";
                when x"1CB3" => data <= "00000";
                when x"1CB4" => data <= "00110";
                when x"1CB5" => data <= "00000";
                when x"1CB6" => data <= "00000";
                when x"1CB7" => data <= "00000";
                when x"1CB8" => data <= "00000";
                when x"1CB9" => data <= "00110";
                when x"1CBA" => data <= "00000";
                when x"1CBB" => data <= "00110";
                when x"1CBC" => data <= "00000";
                when x"1CBD" => data <= "00000";
                when x"1CBE" => data <= "00110";
                when x"1CBF" => data <= "01011";
                when x"1CC0" => data <= "00000";
                when x"1CC1" => data <= "00000";
                when x"1CC2" => data <= "00110";
                when x"1CC3" => data <= "00000";
                when x"1CC4" => data <= "00110";
                when x"1CC5" => data <= "00110";
                when x"1CC6" => data <= "00110";
                when x"1CC7" => data <= "00110";
                when x"1CC8" => data <= "00000";
                when x"1CC9" => data <= "01101";
                when x"1CCA" => data <= "00000";
                when x"1CCB" => data <= "00000";
                when x"1CCC" => data <= "00000";
                when x"1CCD" => data <= "00011";
                when x"1CCE" => data <= "00101";
                when x"1CCF" => data <= "00110";
                when x"1CD0" => data <= "00000";
                when x"1CD1" => data <= "00110";
                when x"1CD2" => data <= "00000";
                when x"1CD3" => data <= "00110";
                when x"1CD4" => data <= "00110";
                when x"1CD5" => data <= "00001";
                when x"1CD6" => data <= "00110";
                when x"1CD7" => data <= "11110";
                when x"1CD8" => data <= "00110";
                when x"1CD9" => data <= "00000";
                when x"1CDA" => data <= "00110";
                when x"1CDB" => data <= "00000";
                when x"1CDC" => data <= "01110";
                when x"1CDD" => data <= "10111";
                when x"1CDE" => data <= "00000";
                when x"1CDF" => data <= "00000";
                when x"1CE0" => data <= "00101";
                when x"1CE1" => data <= "00000";
                when x"1CE2" => data <= "00000";
                when x"1CE3" => data <= "00110";
                when x"1CE4" => data <= "00110";
                when x"1CE5" => data <= "00000";
                when x"1CE6" => data <= "00000";
                when x"1CE7" => data <= "00000";
                when x"1CE8" => data <= "00110";
                when x"1CE9" => data <= "00000";
                when x"1CEA" => data <= "00110";
                when x"1CEB" => data <= "00110";
                when x"1CEC" => data <= "00000";
                when x"1CED" => data <= "10101";
                when x"1CEE" => data <= "11100";
                when x"1CEF" => data <= "00110";
                when x"1CF0" => data <= "00000";
                when x"1CF1" => data <= "00110";
                when x"1CF2" => data <= "00110";
                when x"1CF3" => data <= "00000";
                when x"1CF4" => data <= "00110";
                when x"1CF5" => data <= "00110";
                when x"1CF6" => data <= "00000";
                when x"1CF7" => data <= "00110";
                when x"1CF8" => data <= "00110";
                when x"1CF9" => data <= "00000";
                when x"1CFA" => data <= "00110";
                when x"1CFB" => data <= "01010";
                when x"1CFC" => data <= "00110";
                when x"1CFD" => data <= "00110";
                when x"1CFE" => data <= "01011";
                when x"1CFF" => data <= "01101";
                when x"1D00" => data <= "00110";
                when x"1D01" => data <= "00000";
                when x"1D02" => data <= "00000";
                when x"1D03" => data <= "00110";
                when x"1D04" => data <= "00110";
                when x"1D05" => data <= "00110";
                when x"1D06" => data <= "00110";
                when x"1D07" => data <= "00110";
                when x"1D08" => data <= "00000";
                when x"1D09" => data <= "10100";
                when x"1D0A" => data <= "00110";
                when x"1D0B" => data <= "00000";
                when x"1D0C" => data <= "00000";
                when x"1D0D" => data <= "00110";
                when x"1D0E" => data <= "11001";
                when x"1D0F" => data <= "00111";
                when x"1D10" => data <= "00110";
                when x"1D11" => data <= "00000";
                when x"1D12" => data <= "00000";
                when x"1D13" => data <= "00000";
                when x"1D14" => data <= "01011";
                when x"1D15" => data <= "00110";
                when x"1D16" => data <= "00000";
                when x"1D17" => data <= "00110";
                when x"1D18" => data <= "00110";
                when x"1D19" => data <= "00110";
                when x"1D1A" => data <= "00000";
                when x"1D1B" => data <= "00000";
                when x"1D1C" => data <= "00000";
                when x"1D1D" => data <= "00110";
                when x"1D1E" => data <= "00000";
                when x"1D1F" => data <= "00000";
                when x"1D20" => data <= "00110";
                when x"1D21" => data <= "00110";
                when x"1D22" => data <= "00110";
                when x"1D23" => data <= "00110";
                when x"1D24" => data <= "10000";
                when x"1D25" => data <= "00110";
                when x"1D26" => data <= "01001";
                when x"1D27" => data <= "10011";
                when x"1D28" => data <= "00110";
                when x"1D29" => data <= "00000";
                when x"1D2A" => data <= "00000";
                when x"1D2B" => data <= "00000";
                when x"1D2C" => data <= "00000";
                when x"1D2D" => data <= "00000";
                when x"1D2E" => data <= "00110";
                when x"1D2F" => data <= "00000";
                when x"1D30" => data <= "00110";
                when x"1D31" => data <= "00110";
                when x"1D32" => data <= "00000";
                when x"1D33" => data <= "00000";
                when x"1D34" => data <= "01100";
                when x"1D35" => data <= "00110";
                when x"1D36" => data <= "01011";
                when x"1D37" => data <= "00000";
                when x"1D38" => data <= "00000";
                when x"1D39" => data <= "00000";
                when x"1D3A" => data <= "00110";
                when x"1D3B" => data <= "00000";
                when x"1D3C" => data <= "00000";
                when x"1D3D" => data <= "00110";
                when x"1D3E" => data <= "00110";
                when x"1D3F" => data <= "00000";
                when x"1D40" => data <= "00110";
                when x"1D41" => data <= "00000";
                when x"1D42" => data <= "00110";
                when x"1D43" => data <= "11001";
                when x"1D44" => data <= "00110";
                when x"1D45" => data <= "00011";
                when x"1D46" => data <= "11110";
                when x"1D47" => data <= "00000";
                when x"1D48" => data <= "00000";
                when x"1D49" => data <= "00110";
                when x"1D4A" => data <= "01101";
                when x"1D4B" => data <= "00000";
                when x"1D4C" => data <= "00000";
                when x"1D4D" => data <= "00000";
                when x"1D4E" => data <= "00000";
                when x"1D4F" => data <= "11010";
                when x"1D50" => data <= "00000";
                when x"1D51" => data <= "00110";
                when x"1D52" => data <= "00110";
                when x"1D53" => data <= "00110";
                when x"1D54" => data <= "00110";
                when x"1D55" => data <= "00001";
                when x"1D56" => data <= "00110";
                when x"1D57" => data <= "10000";
                when x"1D58" => data <= "01011";
                when x"1D59" => data <= "00110";
                when x"1D5A" => data <= "00110";
                when x"1D5B" => data <= "00110";
                when x"1D5C" => data <= "10011";
                when x"1D5D" => data <= "00000";
                when x"1D5E" => data <= "00110";
                when x"1D5F" => data <= "00000";
                when x"1D60" => data <= "00000";
                when x"1D61" => data <= "00000";
                when x"1D62" => data <= "00110";
                when x"1D63" => data <= "00110";
                when x"1D64" => data <= "00110";
                when x"1D65" => data <= "00000";
                when x"1D66" => data <= "10011";
                when x"1D67" => data <= "11111";
                when x"1D68" => data <= "00000";
                when x"1D69" => data <= "00110";
                when x"1D6A" => data <= "00000";
                when x"1D6B" => data <= "00000";
                when x"1D6C" => data <= "00110";
                when x"1D6D" => data <= "00110";
                when x"1D6E" => data <= "01110";
                when x"1D6F" => data <= "00000";
                when x"1D70" => data <= "00110";
                when x"1D71" => data <= "00000";
                when x"1D72" => data <= "00110";
                when x"1D73" => data <= "00000";
                when x"1D74" => data <= "01101";
                when x"1D75" => data <= "00000";
                when x"1D76" => data <= "00000";
                when x"1D77" => data <= "00000";
                when x"1D78" => data <= "00110";
                when x"1D79" => data <= "00110";
                when x"1D7A" => data <= "00110";
                when x"1D7B" => data <= "00000";
                when x"1D7C" => data <= "00000";
                when x"1D7D" => data <= "00000";
                when x"1D7E" => data <= "00110";
                when x"1D7F" => data <= "00000";
                when x"1D80" => data <= "00000";
                when x"1D81" => data <= "00110";
                when x"1D82" => data <= "00000";
                when x"1D83" => data <= "00110";
                when x"1D84" => data <= "00110";
                when x"1D85" => data <= "00110";
                when x"1D86" => data <= "01011";
                when x"1D87" => data <= "00110";
                when x"1D88" => data <= "01011";
                when x"1D89" => data <= "00110";
                when x"1D8A" => data <= "00110";
                when x"1D8B" => data <= "00110";
                when x"1D8C" => data <= "00110";
                when x"1D8D" => data <= "00110";
                when x"1D8E" => data <= "00110";
                when x"1D8F" => data <= "01000";
                when x"1D90" => data <= "00110";
                when x"1D91" => data <= "01110";
                when x"1D92" => data <= "01110";
                when x"1D93" => data <= "00000";
                when x"1D94" => data <= "01001";
                when x"1D95" => data <= "00000";
                when x"1D96" => data <= "00110";
                when x"1D97" => data <= "00000";
                when x"1D98" => data <= "00000";
                when x"1D99" => data <= "00000";
                when x"1D9A" => data <= "00000";
                when x"1D9B" => data <= "00000";
                when x"1D9C" => data <= "01110";
                when x"1D9D" => data <= "10101";
                when x"1D9E" => data <= "00110";
                when x"1D9F" => data <= "00110";
                when x"1DA0" => data <= "00000";
                when x"1DA1" => data <= "00110";
                when x"1DA2" => data <= "00000";
                when x"1DA3" => data <= "00000";
                when x"1DA4" => data <= "00110";
                when x"1DA5" => data <= "00000";
                when x"1DA6" => data <= "00110";
                when x"1DA7" => data <= "00110";
                when x"1DA8" => data <= "00000";
                when x"1DA9" => data <= "00000";
                when x"1DAA" => data <= "00000";
                when x"1DAB" => data <= "00000";
                when x"1DAC" => data <= "00110";
                when x"1DAD" => data <= "00000";
                when x"1DAE" => data <= "00000";
                when x"1DAF" => data <= "00000";
                when x"1DB0" => data <= "01101";
                when x"1DB1" => data <= "11000";
                when x"1DB2" => data <= "00000";
                when x"1DB3" => data <= "11110";
                when x"1DB4" => data <= "00110";
                when x"1DB5" => data <= "00110";
                when x"1DB6" => data <= "00000";
                when x"1DB7" => data <= "00000";
                when x"1DB8" => data <= "00110";
                when x"1DB9" => data <= "00000";
                when x"1DBA" => data <= "01101";
                when x"1DBB" => data <= "00110";
                when x"1DBC" => data <= "00000";
                when x"1DBD" => data <= "00000";
                when x"1DBE" => data <= "00000";
                when x"1DBF" => data <= "00000";
                when x"1DC0" => data <= "00110";
                when x"1DC1" => data <= "01001";
                when x"1DC2" => data <= "00110";
                when x"1DC3" => data <= "00110";
                when x"1DC4" => data <= "01011";
                when x"1DC5" => data <= "00000";
                when x"1DC6" => data <= "00000";
                when x"1DC7" => data <= "00000";
                when x"1DC8" => data <= "00000";
                when x"1DC9" => data <= "00000";
                when x"1DCA" => data <= "00000";
                when x"1DCB" => data <= "00110";
                when x"1DCC" => data <= "00110";
                when x"1DCD" => data <= "00110";
                when x"1DCE" => data <= "10010";
                when x"1DCF" => data <= "00110";
                when x"1DD0" => data <= "00110";
                when x"1DD1" => data <= "01011";
                when x"1DD2" => data <= "00110";
                when x"1DD3" => data <= "00110";
                when x"1DD4" => data <= "00110";
                when x"1DD5" => data <= "00110";
                when x"1DD6" => data <= "01101";
                when x"1DD7" => data <= "01011";
                when x"1DD8" => data <= "00110";
                when x"1DD9" => data <= "00110";
                when x"1DDA" => data <= "00110";
                when x"1DDB" => data <= "00000";
                when x"1DDC" => data <= "00000";
                when x"1DDD" => data <= "10110";
                when x"1DDE" => data <= "00000";
                when x"1DDF" => data <= "00000";
                when x"1DE0" => data <= "00000";
                when x"1DE1" => data <= "00110";
                when x"1DE2" => data <= "10100";
                when x"1DE3" => data <= "00110";
                when x"1DE4" => data <= "00110";
                when x"1DE5" => data <= "00110";
                when x"1DE6" => data <= "00000";
                when x"1DE7" => data <= "00110";
                when x"1DE8" => data <= "11011";
                when x"1DE9" => data <= "10011";
                when x"1DEA" => data <= "00110";
                when x"1DEB" => data <= "00110";
                when x"1DEC" => data <= "11111";
                when x"1DED" => data <= "00000";
                when x"1DEE" => data <= "00110";
                when x"1DEF" => data <= "10110";
                when x"1DF0" => data <= "00110";
                when x"1DF1" => data <= "00110";
                when x"1DF2" => data <= "00000";
                when x"1DF3" => data <= "01001";
                when x"1DF4" => data <= "00110";
                when x"1DF5" => data <= "00101";
                when x"1DF6" => data <= "00110";
                when x"1DF7" => data <= "00110";
                when x"1DF8" => data <= "00000";
                when x"1DF9" => data <= "00110";
                when x"1DFA" => data <= "00110";
                when x"1DFB" => data <= "00110";
                when x"1DFC" => data <= "11100";
                when x"1DFD" => data <= "00000";
                when x"1DFE" => data <= "00000";
                when x"1DFF" => data <= "00000";
                when x"1E00" => data <= "00000";
                when x"1E01" => data <= "00000";
                when x"1E02" => data <= "00110";
                when x"1E03" => data <= "01011";
                when x"1E04" => data <= "00110";
                when x"1E05" => data <= "11010";
                when x"1E06" => data <= "00000";
                when x"1E07" => data <= "00110";
                when x"1E08" => data <= "00000";
                when x"1E09" => data <= "00110";
                when x"1E0A" => data <= "00000";
                when x"1E0B" => data <= "00110";
                when x"1E0C" => data <= "11101";
                when x"1E0D" => data <= "00000";
                when x"1E0E" => data <= "00000";
                when x"1E0F" => data <= "00000";
                when x"1E10" => data <= "00110";
                when x"1E11" => data <= "00110";
                when x"1E12" => data <= "00000";
                when x"1E13" => data <= "00000";
                when x"1E14" => data <= "01000";
                when x"1E15" => data <= "00000";
                when x"1E16" => data <= "11111";
                when x"1E17" => data <= "00110";
                when x"1E18" => data <= "00000";
                when x"1E19" => data <= "00000";
                when x"1E1A" => data <= "00000";
                when x"1E1B" => data <= "00000";
                when x"1E1C" => data <= "11110";
                when x"1E1D" => data <= "00100";
                when x"1E1E" => data <= "01011";
                when x"1E1F" => data <= "01011";
                when x"1E20" => data <= "10001";
                when x"1E21" => data <= "00110";
                when x"1E22" => data <= "00000";
                when x"1E23" => data <= "00110";
                when x"1E24" => data <= "01010";
                when x"1E25" => data <= "00000";
                when x"1E26" => data <= "00111";
                when x"1E27" => data <= "00110";
                when x"1E28" => data <= "00110";
                when x"1E29" => data <= "00000";
                when x"1E2A" => data <= "00110";
                when x"1E2B" => data <= "00101";
                when x"1E2C" => data <= "00000";
                when x"1E2D" => data <= "00110";
                when x"1E2E" => data <= "00000";
                when x"1E2F" => data <= "00000";
                when x"1E30" => data <= "00000";
                when x"1E31" => data <= "00110";
                when x"1E32" => data <= "00000";
                when x"1E33" => data <= "00110";
                when x"1E34" => data <= "01100";
                when x"1E35" => data <= "00110";
                when x"1E36" => data <= "11000";
                when x"1E37" => data <= "00110";
                when x"1E38" => data <= "01101";
                when x"1E39" => data <= "00000";
                when x"1E3A" => data <= "00110";
                when x"1E3B" => data <= "00000";
                when x"1E3C" => data <= "00000";
                when x"1E3D" => data <= "00110";
                when x"1E3E" => data <= "00110";
                when x"1E3F" => data <= "00000";
                when x"1E40" => data <= "00000";
                when x"1E41" => data <= "00110";
                when x"1E42" => data <= "00000";
                when x"1E43" => data <= "11010";
                when x"1E44" => data <= "00110";
                when x"1E45" => data <= "00000";
                when x"1E46" => data <= "10100";
                when x"1E47" => data <= "11110";
                when x"1E48" => data <= "01011";
                when x"1E49" => data <= "00110";
                when x"1E4A" => data <= "01010";
                when x"1E4B" => data <= "00110";
                when x"1E4C" => data <= "00110";
                when x"1E4D" => data <= "00110";
                when x"1E4E" => data <= "10000";
                when x"1E4F" => data <= "00000";
                when x"1E50" => data <= "00000";
                when x"1E51" => data <= "00110";
                when x"1E52" => data <= "00000";
                when x"1E53" => data <= "00110";
                when x"1E54" => data <= "00000";
                when x"1E55" => data <= "00110";
                when x"1E56" => data <= "00110";
                when x"1E57" => data <= "00110";
                when x"1E58" => data <= "00110";
                when x"1E59" => data <= "00000";
                when x"1E5A" => data <= "00110";
                when x"1E5B" => data <= "00000";
                when x"1E5C" => data <= "00110";
                when x"1E5D" => data <= "11100";
                when x"1E5E" => data <= "00000";
                when x"1E5F" => data <= "00000";
                when x"1E60" => data <= "00110";
                when x"1E61" => data <= "00000";
                when x"1E62" => data <= "00000";
                when x"1E63" => data <= "00000";
                when x"1E64" => data <= "00110";
                when x"1E65" => data <= "00000";
                when x"1E66" => data <= "00000";
                when x"1E67" => data <= "11001";
                when x"1E68" => data <= "00000";
                when x"1E69" => data <= "00110";
                when x"1E6A" => data <= "10011";
                when x"1E6B" => data <= "00110";
                when x"1E6C" => data <= "00110";
                when x"1E6D" => data <= "00110";
                when x"1E6E" => data <= "00110";
                when x"1E6F" => data <= "00110";
                when x"1E70" => data <= "00000";
                when x"1E71" => data <= "00000";
                when x"1E72" => data <= "11000";
                when x"1E73" => data <= "11001";
                when x"1E74" => data <= "00110";
                when x"1E75" => data <= "11111";
                when x"1E76" => data <= "00000";
                when x"1E77" => data <= "11100";
                when x"1E78" => data <= "00000";
                when x"1E79" => data <= "01110";
                when x"1E7A" => data <= "00110";
                when x"1E7B" => data <= "00000";
                when x"1E7C" => data <= "00000";
                when x"1E7D" => data <= "00110";
                when x"1E7E" => data <= "00110";
                when x"1E7F" => data <= "00110";
                when x"1E80" => data <= "00000";
                when x"1E81" => data <= "00000";
                when x"1E82" => data <= "00000";
                when x"1E83" => data <= "01010";
                when x"1E84" => data <= "00110";
                when x"1E85" => data <= "00110";
                when x"1E86" => data <= "00000";
                when x"1E87" => data <= "00000";
                when x"1E88" => data <= "00110";
                when x"1E89" => data <= "00110";
                when x"1E8A" => data <= "10101";
                when x"1E8B" => data <= "00000";
                when x"1E8C" => data <= "00110";
                when x"1E8D" => data <= "00110";
                when x"1E8E" => data <= "00110";
                when x"1E8F" => data <= "00000";
                when x"1E90" => data <= "00000";
                when x"1E91" => data <= "00000";
                when x"1E92" => data <= "00000";
                when x"1E93" => data <= "00000";
                when x"1E94" => data <= "00110";
                when x"1E95" => data <= "01101";
                when x"1E96" => data <= "00110";
                when x"1E97" => data <= "11111";
                when x"1E98" => data <= "00101";
                when x"1E99" => data <= "00000";
                when x"1E9A" => data <= "01011";
                when x"1E9B" => data <= "00000";
                when x"1E9C" => data <= "00000";
                when x"1E9D" => data <= "11110";
                when x"1E9E" => data <= "00000";
                when x"1E9F" => data <= "00110";
                when x"1EA0" => data <= "00001";
                when x"1EA1" => data <= "00110";
                when x"1EA2" => data <= "00110";
                when x"1EA3" => data <= "00110";
                when x"1EA4" => data <= "01110";
                when x"1EA5" => data <= "00110";
                when x"1EA6" => data <= "10001";
                when x"1EA7" => data <= "00110";
                when x"1EA8" => data <= "10010";
                when x"1EA9" => data <= "00000";
                when x"1EAA" => data <= "00000";
                when x"1EAB" => data <= "00000";
                when x"1EAC" => data <= "00000";
                when x"1EAD" => data <= "00110";
                when x"1EAE" => data <= "00000";
                when x"1EAF" => data <= "00000";
                when x"1EB0" => data <= "00110";
                when x"1EB1" => data <= "00110";
                when x"1EB2" => data <= "10110";
                when x"1EB3" => data <= "00000";
                when x"1EB4" => data <= "00000";
                when x"1EB5" => data <= "00110";
                when x"1EB6" => data <= "00000";
                when x"1EB7" => data <= "00110";
                when x"1EB8" => data <= "00000";
                when x"1EB9" => data <= "10111";
                when x"1EBA" => data <= "00110";
                when x"1EBB" => data <= "00110";
                when x"1EBC" => data <= "01001";
                when x"1EBD" => data <= "00000";
                when x"1EBE" => data <= "00000";
                when x"1EBF" => data <= "00110";
                when x"1EC0" => data <= "00000";
                when x"1EC1" => data <= "01101";
                when x"1EC2" => data <= "00000";
                when x"1EC3" => data <= "00000";
                when x"1EC4" => data <= "00110";
                when x"1EC5" => data <= "00110";
                when x"1EC6" => data <= "00110";
                when x"1EC7" => data <= "00000";
                when x"1EC8" => data <= "00000";
                when x"1EC9" => data <= "00000";
                when x"1ECA" => data <= "00000";
                when x"1ECB" => data <= "00000";
                when x"1ECC" => data <= "00000";
                when x"1ECD" => data <= "00110";
                when x"1ECE" => data <= "00000";
                when x"1ECF" => data <= "00110";
                when x"1ED0" => data <= "11010";
                when x"1ED1" => data <= "00000";
                when x"1ED2" => data <= "00010";
                when x"1ED3" => data <= "01101";
                when x"1ED4" => data <= "00110";
                when x"1ED5" => data <= "00000";
                when x"1ED6" => data <= "00000";
                when x"1ED7" => data <= "01101";
                when x"1ED8" => data <= "01110";
                when x"1ED9" => data <= "00000";
                when x"1EDA" => data <= "00000";
                when x"1EDB" => data <= "01101";
                when x"1EDC" => data <= "00000";
                when x"1EDD" => data <= "00110";
                when x"1EDE" => data <= "00110";
                when x"1EDF" => data <= "00110";
                when x"1EE0" => data <= "01101";
                when x"1EE1" => data <= "10011";
                when x"1EE2" => data <= "00110";
                when x"1EE3" => data <= "00000";
                when x"1EE4" => data <= "00000";
                when x"1EE5" => data <= "00000";
                when x"1EE6" => data <= "00000";
                when x"1EE7" => data <= "11110";
                when x"1EE8" => data <= "10100";
                when x"1EE9" => data <= "00110";
                when x"1EEA" => data <= "11000";
                when x"1EEB" => data <= "11000";
                when x"1EEC" => data <= "00110";
                when x"1EED" => data <= "00000";
                when x"1EEE" => data <= "00000";
                when x"1EEF" => data <= "00110";
                when x"1EF0" => data <= "01011";
                when x"1EF1" => data <= "00110";
                when x"1EF2" => data <= "00000";
                when x"1EF3" => data <= "10111";
                when x"1EF4" => data <= "00000";
                when x"1EF5" => data <= "00110";
                when x"1EF6" => data <= "00000";
                when x"1EF7" => data <= "00000";
                when x"1EF8" => data <= "00110";
                when x"1EF9" => data <= "00110";
                when x"1EFA" => data <= "00110";
                when x"1EFB" => data <= "10111";
                when x"1EFC" => data <= "01101";
                when x"1EFD" => data <= "01011";
                when x"1EFE" => data <= "00110";
                when x"1EFF" => data <= "00110";
                when x"1F00" => data <= "01011";
                when x"1F01" => data <= "00000";
                when x"1F02" => data <= "00101";
                when x"1F03" => data <= "00000";
                when x"1F04" => data <= "01001";
                when x"1F05" => data <= "11001";
                when x"1F06" => data <= "00110";
                when x"1F07" => data <= "00110";
                when x"1F08" => data <= "01010";
                when x"1F09" => data <= "00000";
                when x"1F0A" => data <= "00110";
                when x"1F0B" => data <= "00011";
                when x"1F0C" => data <= "00000";
                when x"1F0D" => data <= "00110";
                when x"1F0E" => data <= "10100";
                when x"1F0F" => data <= "00110";
                when x"1F10" => data <= "00000";
                when x"1F11" => data <= "00000";
                when x"1F12" => data <= "11010";
                when x"1F13" => data <= "00110";
                when x"1F14" => data <= "00110";
                when x"1F15" => data <= "00110";
                when x"1F16" => data <= "01100";
                when x"1F17" => data <= "00110";
                when x"1F18" => data <= "00000";
                when x"1F19" => data <= "00000";
                when x"1F1A" => data <= "00110";
                when x"1F1B" => data <= "00000";
                when x"1F1C" => data <= "00000";
                when x"1F1D" => data <= "00110";
                when x"1F1E" => data <= "00110";
                when x"1F1F" => data <= "00100";
                when x"1F20" => data <= "00110";
                when x"1F21" => data <= "00000";
                when x"1F22" => data <= "00000";
                when x"1F23" => data <= "00000";
                when x"1F24" => data <= "00101";
                when x"1F25" => data <= "00110";
                when x"1F26" => data <= "01000";
                when x"1F27" => data <= "00110";
                when x"1F28" => data <= "10011";
                when x"1F29" => data <= "00000";
                when x"1F2A" => data <= "00110";
                when x"1F2B" => data <= "00110";
                when x"1F2C" => data <= "00000";
                when x"1F2D" => data <= "00110";
                when x"1F2E" => data <= "00110";
                when x"1F2F" => data <= "00000";
                when x"1F30" => data <= "00000";
                when x"1F31" => data <= "00110";
                when x"1F32" => data <= "00000";
                when x"1F33" => data <= "10010";
                when x"1F34" => data <= "00110";
                when x"1F35" => data <= "00000";
                when x"1F36" => data <= "00110";
                when x"1F37" => data <= "00110";
                when x"1F38" => data <= "00110";
                when x"1F39" => data <= "00000";
                when x"1F3A" => data <= "00000";
                when x"1F3B" => data <= "00000";
                when x"1F3C" => data <= "00000";
                when x"1F3D" => data <= "00000";
                when x"1F3E" => data <= "00000";
                when x"1F3F" => data <= "00110";
                when x"1F40" => data <= "00110";
                when x"1F41" => data <= "01101";
                when x"1F42" => data <= "00000";
                when x"1F43" => data <= "00110";
                when x"1F44" => data <= "01100";
                when x"1F45" => data <= "00000";
                when x"1F46" => data <= "00110";
                when x"1F47" => data <= "00110";
                when x"1F48" => data <= "00000";
                when x"1F49" => data <= "11001";
                when x"1F4A" => data <= "00000";
                when x"1F4B" => data <= "00110";
                when x"1F4C" => data <= "00000";
                when x"1F4D" => data <= "01101";
                when x"1F4E" => data <= "00000";
                when x"1F4F" => data <= "11110";
                when x"1F50" => data <= "00110";
                when x"1F51" => data <= "00110";
                when x"1F52" => data <= "00110";
                when x"1F53" => data <= "00000";
                when x"1F54" => data <= "00110";
                when x"1F55" => data <= "00110";
                when x"1F56" => data <= "00000";
                when x"1F57" => data <= "00110";
                when x"1F58" => data <= "00110";
                when x"1F59" => data <= "10001";
                when x"1F5A" => data <= "00110";
                when x"1F5B" => data <= "00110";
                when x"1F5C" => data <= "00110";
                when x"1F5D" => data <= "00110";
                when x"1F5E" => data <= "00110";
                when x"1F5F" => data <= "00000";
                when x"1F60" => data <= "00110";
                when x"1F61" => data <= "00000";
                when x"1F62" => data <= "10001";
                when x"1F63" => data <= "00000";
                when x"1F64" => data <= "00000";
                when x"1F65" => data <= "00110";
                when x"1F66" => data <= "00000";
                when x"1F67" => data <= "00000";
                when x"1F68" => data <= "00110";
                when x"1F69" => data <= "00110";
                when x"1F6A" => data <= "00000";
                when x"1F6B" => data <= "00000";
                when x"1F6C" => data <= "00000";
                when x"1F6D" => data <= "00000";
                when x"1F6E" => data <= "00000";
                when x"1F6F" => data <= "00110";
                when x"1F70" => data <= "00110";
                when x"1F71" => data <= "00110";
                when x"1F72" => data <= "00110";
                when x"1F73" => data <= "00000";
                when x"1F74" => data <= "00000";
                when x"1F75" => data <= "00110";
                when x"1F76" => data <= "00000";
                when x"1F77" => data <= "00000";
                when x"1F78" => data <= "00000";
                when x"1F79" => data <= "11110";
                when x"1F7A" => data <= "10010";
                when x"1F7B" => data <= "00000";
                when x"1F7C" => data <= "00000";
                when x"1F7D" => data <= "00110";
                when x"1F7E" => data <= "00000";
                when x"1F7F" => data <= "11001";
                when x"1F80" => data <= "00000";
                when x"1F81" => data <= "00110";
                when x"1F82" => data <= "00000";
                when x"1F83" => data <= "00000";
                when x"1F84" => data <= "00000";
                when x"1F85" => data <= "00110";
                when x"1F86" => data <= "00000";
                when x"1F87" => data <= "00110";
                when x"1F88" => data <= "00000";
                when x"1F89" => data <= "01001";
                when x"1F8A" => data <= "10101";
                when x"1F8B" => data <= "00110";
                when x"1F8C" => data <= "00110";
                when x"1F8D" => data <= "00110";
                when x"1F8E" => data <= "00000";
                when x"1F8F" => data <= "00000";
                when x"1F90" => data <= "00110";
                when x"1F91" => data <= "00000";
                when x"1F92" => data <= "00000";
                when x"1F93" => data <= "00110";
                when x"1F94" => data <= "00000";
                when x"1F95" => data <= "00000";
                when x"1F96" => data <= "00110";
                when x"1F97" => data <= "00000";
                when x"1F98" => data <= "00110";
                when x"1F99" => data <= "00110";
                when x"1F9A" => data <= "00010";
                when x"1F9B" => data <= "11100";
                when x"1F9C" => data <= "01110";
                when x"1F9D" => data <= "00000";
                when x"1F9E" => data <= "10011";
                when x"1F9F" => data <= "00000";
                when x"1FA0" => data <= "00000";
                when x"1FA1" => data <= "00000";
                when x"1FA2" => data <= "10101";
                when x"1FA3" => data <= "00110";
                when x"1FA4" => data <= "00101";
                when x"1FA5" => data <= "01111";
                when x"1FA6" => data <= "00000";
                when x"1FA7" => data <= "00110";
                when x"1FA8" => data <= "10000";
                when x"1FA9" => data <= "00101";
                when x"1FAA" => data <= "00110";
                when x"1FAB" => data <= "11110";
                when x"1FAC" => data <= "00110";
                when x"1FAD" => data <= "00110";
                when x"1FAE" => data <= "00110";
                when x"1FAF" => data <= "00110";
                when x"1FB0" => data <= "00110";
                when x"1FB1" => data <= "01011";
                when x"1FB2" => data <= "00110";
                when x"1FB3" => data <= "00000";
                when x"1FB4" => data <= "00001";
                when x"1FB5" => data <= "00110";
                when x"1FB6" => data <= "01000";
                when x"1FB7" => data <= "01010";
                when x"1FB8" => data <= "00110";
                when x"1FB9" => data <= "00110";
                when x"1FBA" => data <= "10110";
                when x"1FBB" => data <= "00110";
                when x"1FBC" => data <= "00000";
                when x"1FBD" => data <= "00110";
                when x"1FBE" => data <= "00110";
                when x"1FBF" => data <= "00000";
                when x"1FC0" => data <= "00110";
                when x"1FC1" => data <= "00110";
                when x"1FC2" => data <= "00000";
                when x"1FC3" => data <= "00110";
                when x"1FC4" => data <= "00000";
                when x"1FC5" => data <= "00110";
                when x"1FC6" => data <= "00110";
                when x"1FC7" => data <= "00110";
                when x"1FC8" => data <= "00110";
                when x"1FC9" => data <= "00110";
                when x"1FCA" => data <= "10111";
                when x"1FCB" => data <= "00000";
                when x"1FCC" => data <= "00000";
                when x"1FCD" => data <= "00000";
                when x"1FCE" => data <= "00000";
                when x"1FCF" => data <= "00000";
                when x"1FD0" => data <= "00000";
                when x"1FD1" => data <= "10101";
                when x"1FD2" => data <= "11001";
                when x"1FD3" => data <= "01000";
                when x"1FD4" => data <= "00000";
                when x"1FD5" => data <= "00000";
                when x"1FD6" => data <= "00000";
                when x"1FD7" => data <= "00110";
                when x"1FD8" => data <= "00110";
                when x"1FD9" => data <= "00110";
                when x"1FDA" => data <= "01010";
                when x"1FDB" => data <= "00110";
                when x"1FDC" => data <= "00110";
                when x"1FDD" => data <= "01111";
                when x"1FDE" => data <= "00000";
                when x"1FDF" => data <= "00000";
                when x"1FE0" => data <= "00110";
                when x"1FE1" => data <= "00110";
                when x"1FE2" => data <= "00110";
                when x"1FE3" => data <= "00110";
                when x"1FE4" => data <= "00000";
                when x"1FE5" => data <= "01110";
                when x"1FE6" => data <= "00000";
                when x"1FE7" => data <= "00000";
                when x"1FE8" => data <= "00110";
                when x"1FE9" => data <= "00000";
                when x"1FEA" => data <= "00110";
                when x"1FEB" => data <= "00001";
                when x"1FEC" => data <= "00000";
                when x"1FED" => data <= "00011";
                when x"1FEE" => data <= "01111";
                when x"1FEF" => data <= "00110";
                when x"1FF0" => data <= "00110";
                when x"1FF1" => data <= "00110";
                when x"1FF2" => data <= "00000";
                when x"1FF3" => data <= "00000";
                when x"1FF4" => data <= "00000";
                when x"1FF5" => data <= "00110";
                when x"1FF6" => data <= "00000";
                when x"1FF7" => data <= "00110";
                when x"1FF8" => data <= "00110";
                when x"1FF9" => data <= "00110";
                when x"1FFA" => data <= "11111";
                when x"1FFB" => data <= "00110";
                when x"1FFC" => data <= "00000";
                when x"1FFD" => data <= "00110";
                when x"1FFE" => data <= "11100";
                when x"1FFF" => data <= "01101";
                when x"2000" => data <= "00110";
                when x"2001" => data <= "00011";
                when x"2002" => data <= "00000";
                when x"2003" => data <= "01100";
                when x"2004" => data <= "00000";
                when x"2005" => data <= "00011";
                when x"2006" => data <= "01011";
                when x"2007" => data <= "00000";
                when x"2008" => data <= "01101";
                when x"2009" => data <= "00000";
                when x"200A" => data <= "00110";
                when x"200B" => data <= "00110";
                when x"200C" => data <= "00111";
                when x"200D" => data <= "00110";
                when x"200E" => data <= "01010";
                when x"200F" => data <= "11001";
                when x"2010" => data <= "00000";
                when x"2011" => data <= "00000";
                when x"2012" => data <= "00110";
                when x"2013" => data <= "00000";
                when x"2014" => data <= "00110";
                when x"2015" => data <= "11110";
                when x"2016" => data <= "00000";
                when x"2017" => data <= "00000";
                when x"2018" => data <= "00000";
                when x"2019" => data <= "00110";
                when x"201A" => data <= "00110";
                when x"201B" => data <= "01101";
                when x"201C" => data <= "00000";
                when x"201D" => data <= "00110";
                when x"201E" => data <= "01000";
                when x"201F" => data <= "00110";
                when x"2020" => data <= "00000";
                when x"2021" => data <= "00000";
                when x"2022" => data <= "00110";
                when x"2023" => data <= "00000";
                when x"2024" => data <= "01101";
                when x"2025" => data <= "00000";
                when x"2026" => data <= "11011";
                when x"2027" => data <= "01011";
                when x"2028" => data <= "00000";
                when x"2029" => data <= "00110";
                when x"202A" => data <= "01011";
                when x"202B" => data <= "10011";
                when x"202C" => data <= "00000";
                when x"202D" => data <= "00011";
                when x"202E" => data <= "01011";
                when x"202F" => data <= "00000";
                when x"2030" => data <= "00000";
                when x"2031" => data <= "00110";
                when x"2032" => data <= "10010";
                when x"2033" => data <= "00110";
                when x"2034" => data <= "00110";
                when x"2035" => data <= "00110";
                when x"2036" => data <= "00000";
                when x"2037" => data <= "00000";
                when x"2038" => data <= "00000";
                when x"2039" => data <= "00000";
                when x"203A" => data <= "00000";
                when x"203B" => data <= "00110";
                when x"203C" => data <= "00111";
                when x"203D" => data <= "00110";
                when x"203E" => data <= "00000";
                when x"203F" => data <= "00110";
                when x"2040" => data <= "00110";
                when x"2041" => data <= "01000";
                when x"2042" => data <= "10000";
                when x"2043" => data <= "10001";
                when x"2044" => data <= "00000";
                when x"2045" => data <= "00000";
                when x"2046" => data <= "00110";
                when x"2047" => data <= "00111";
                when x"2048" => data <= "00000";
                when x"2049" => data <= "00000";
                when x"204A" => data <= "01101";
                when x"204B" => data <= "01100";
                when x"204C" => data <= "00110";
                when x"204D" => data <= "00000";
                when x"204E" => data <= "00110";
                when x"204F" => data <= "00110";
                when x"2050" => data <= "00000";
                when x"2051" => data <= "10110";
                when x"2052" => data <= "00000";
                when x"2053" => data <= "00000";
                when x"2054" => data <= "00000";
                when x"2055" => data <= "00110";
                when x"2056" => data <= "00110";
                when x"2057" => data <= "00110";
                when x"2058" => data <= "00000";
                when x"2059" => data <= "00110";
                when x"205A" => data <= "10110";
                when x"205B" => data <= "00111";
                when x"205C" => data <= "00000";
                when x"205D" => data <= "00110";
                when x"205E" => data <= "00101";
                when x"205F" => data <= "01011";
                when x"2060" => data <= "00110";
                when x"2061" => data <= "00000";
                when x"2062" => data <= "00000";
                when x"2063" => data <= "00000";
                when x"2064" => data <= "00000";
                when x"2065" => data <= "00000";
                when x"2066" => data <= "10110";
                when x"2067" => data <= "00000";
                when x"2068" => data <= "00000";
                when x"2069" => data <= "00110";
                when x"206A" => data <= "11000";
                when x"206B" => data <= "00110";
                when x"206C" => data <= "00110";
                when x"206D" => data <= "00110";
                when x"206E" => data <= "00110";
                when x"206F" => data <= "00001";
                when x"2070" => data <= "00110";
                when x"2071" => data <= "00000";
                when x"2072" => data <= "00110";
                when x"2073" => data <= "00110";
                when x"2074" => data <= "01101";
                when x"2075" => data <= "10000";
                when x"2076" => data <= "00000";
                when x"2077" => data <= "01111";
                when x"2078" => data <= "00110";
                when x"2079" => data <= "00110";
                when x"207A" => data <= "00110";
                when x"207B" => data <= "00110";
                when x"207C" => data <= "00110";
                when x"207D" => data <= "00000";
                when x"207E" => data <= "00110";
                when x"207F" => data <= "00000";
                when x"2080" => data <= "00000";
                when x"2081" => data <= "01110";
                when x"2082" => data <= "00110";
                when x"2083" => data <= "00000";
                when x"2084" => data <= "01011";
                when x"2085" => data <= "00001";
                when x"2086" => data <= "00000";
                when x"2087" => data <= "00110";
                when x"2088" => data <= "00110";
                when x"2089" => data <= "00000";
                when x"208A" => data <= "00000";
                when x"208B" => data <= "00000";
                when x"208C" => data <= "00110";
                when x"208D" => data <= "00000";
                when x"208E" => data <= "00000";
                when x"208F" => data <= "00110";
                when x"2090" => data <= "00000";
                when x"2091" => data <= "00110";
                when x"2092" => data <= "00110";
                when x"2093" => data <= "10001";
                when x"2094" => data <= "00000";
                when x"2095" => data <= "00000";
                when x"2096" => data <= "00000";
                when x"2097" => data <= "00000";
                when x"2098" => data <= "01100";
                when x"2099" => data <= "00000";
                when x"209A" => data <= "01100";
                when x"209B" => data <= "00000";
                when x"209C" => data <= "00001";
                when x"209D" => data <= "00110";
                when x"209E" => data <= "00110";
                when x"209F" => data <= "00110";
                when x"20A0" => data <= "00110";
                when x"20A1" => data <= "00000";
                when x"20A2" => data <= "00110";
                when x"20A3" => data <= "00000";
                when x"20A4" => data <= "00000";
                when x"20A5" => data <= "00110";
                when x"20A6" => data <= "00110";
                when x"20A7" => data <= "11000";
                when x"20A8" => data <= "11001";
                when x"20A9" => data <= "00000";
                when x"20AA" => data <= "10001";
                when x"20AB" => data <= "00110";
                when x"20AC" => data <= "00000";
                when x"20AD" => data <= "01011";
                when x"20AE" => data <= "00110";
                when x"20AF" => data <= "00000";
                when x"20B0" => data <= "00000";
                when x"20B1" => data <= "00110";
                when x"20B2" => data <= "00110";
                when x"20B3" => data <= "00110";
                when x"20B4" => data <= "01110";
                when x"20B5" => data <= "01000";
                when x"20B6" => data <= "00110";
                when x"20B7" => data <= "00000";
                when x"20B8" => data <= "00000";
                when x"20B9" => data <= "00000";
                when x"20BA" => data <= "01111";
                when x"20BB" => data <= "00110";
                when x"20BC" => data <= "00110";
                when x"20BD" => data <= "00000";
                when x"20BE" => data <= "00000";
                when x"20BF" => data <= "00110";
                when x"20C0" => data <= "00110";
                when x"20C1" => data <= "00110";
                when x"20C2" => data <= "00110";
                when x"20C3" => data <= "00110";
                when x"20C4" => data <= "00000";
                when x"20C5" => data <= "00110";
                when x"20C6" => data <= "00110";
                when x"20C7" => data <= "01001";
                when x"20C8" => data <= "00000";
                when x"20C9" => data <= "00110";
                when x"20CA" => data <= "00000";
                when x"20CB" => data <= "10010";
                when x"20CC" => data <= "01011";
                when x"20CD" => data <= "00110";
                when x"20CE" => data <= "00101";
                when x"20CF" => data <= "01111";
                when x"20D0" => data <= "00000";
                when x"20D1" => data <= "00110";
                when x"20D2" => data <= "00000";
                when x"20D3" => data <= "00000";
                when x"20D4" => data <= "00110";
                when x"20D5" => data <= "01111";
                when x"20D6" => data <= "00000";
                when x"20D7" => data <= "00000";
                when x"20D8" => data <= "00000";
                when x"20D9" => data <= "00000";
                when x"20DA" => data <= "00111";
                when x"20DB" => data <= "00110";
                when x"20DC" => data <= "00000";
                when x"20DD" => data <= "00000";
                when x"20DE" => data <= "00110";
                when x"20DF" => data <= "00110";
                when x"20E0" => data <= "00110";
                when x"20E1" => data <= "00000";
                when x"20E2" => data <= "11101";
                when x"20E3" => data <= "00110";
                when x"20E4" => data <= "00000";
                when x"20E5" => data <= "00000";
                when x"20E6" => data <= "00000";
                when x"20E7" => data <= "01010";
                when x"20E8" => data <= "00110";
                when x"20E9" => data <= "00000";
                when x"20EA" => data <= "00110";
                when x"20EB" => data <= "00100";
                when x"20EC" => data <= "00000";
                when x"20ED" => data <= "00110";
                when x"20EE" => data <= "00000";
                when x"20EF" => data <= "00000";
                when x"20F0" => data <= "00110";
                when x"20F1" => data <= "00000";
                when x"20F2" => data <= "00010";
                when x"20F3" => data <= "00110";
                when x"20F4" => data <= "11111";
                when x"20F5" => data <= "00000";
                when x"20F6" => data <= "11111";
                when x"20F7" => data <= "00000";
                when x"20F8" => data <= "00000";
                when x"20F9" => data <= "00000";
                when x"20FA" => data <= "11110";
                when x"20FB" => data <= "00000";
                when x"20FC" => data <= "00000";
                when x"20FD" => data <= "11000";
                when x"20FE" => data <= "00000";
                when x"20FF" => data <= "00110";
                when x"2100" => data <= "10010";
                when x"2101" => data <= "00110";
                when x"2102" => data <= "00000";
                when x"2103" => data <= "00110";
                when x"2104" => data <= "00000";
                when x"2105" => data <= "00000";
                when x"2106" => data <= "11111";
                when x"2107" => data <= "01100";
                when x"2108" => data <= "00110";
                when x"2109" => data <= "00000";
                when x"210A" => data <= "00000";
                when x"210B" => data <= "00000";
                when x"210C" => data <= "00000";
                when x"210D" => data <= "01011";
                when x"210E" => data <= "00000";
                when x"210F" => data <= "11000";
                when x"2110" => data <= "11001";
                when x"2111" => data <= "00110";
                when x"2112" => data <= "00110";
                when x"2113" => data <= "11111";
                when x"2114" => data <= "00000";
                when x"2115" => data <= "00000";
                when x"2116" => data <= "00000";
                when x"2117" => data <= "00000";
                when x"2118" => data <= "00110";
                when x"2119" => data <= "00000";
                when x"211A" => data <= "00110";
                when x"211B" => data <= "11101";
                when x"211C" => data <= "00000";
                when x"211D" => data <= "00000";
                when x"211E" => data <= "01101";
                when x"211F" => data <= "00000";
                when x"2120" => data <= "00110";
                when x"2121" => data <= "00001";
                when x"2122" => data <= "00000";
                when x"2123" => data <= "11000";
                when x"2124" => data <= "00000";
                when x"2125" => data <= "01000";
                when x"2126" => data <= "11100";
                when x"2127" => data <= "00000";
                when x"2128" => data <= "10011";
                when x"2129" => data <= "00110";
                when x"212A" => data <= "10110";
                when x"212B" => data <= "00000";
                when x"212C" => data <= "00110";
                when x"212D" => data <= "00000";
                when x"212E" => data <= "01111";
                when x"212F" => data <= "00000";
                when x"2130" => data <= "00110";
                when x"2131" => data <= "00110";
                when x"2132" => data <= "11111";
                when x"2133" => data <= "00110";
                when x"2134" => data <= "00000";
                when x"2135" => data <= "00000";
                when x"2136" => data <= "00110";
                when x"2137" => data <= "01010";
                when x"2138" => data <= "00000";
                when x"2139" => data <= "00000";
                when x"213A" => data <= "00000";
                when x"213B" => data <= "10010";
                when x"213C" => data <= "11000";
                when x"213D" => data <= "00000";
                when x"213E" => data <= "00110";
                when x"213F" => data <= "11011";
                when x"2140" => data <= "00000";
                when x"2141" => data <= "00110";
                when x"2142" => data <= "01001";
                when x"2143" => data <= "00110";
                when x"2144" => data <= "00000";
                when x"2145" => data <= "00110";
                when x"2146" => data <= "00110";
                when x"2147" => data <= "00000";
                when x"2148" => data <= "00110";
                when x"2149" => data <= "00110";
                when x"214A" => data <= "00110";
                when x"214B" => data <= "00000";
                when x"214C" => data <= "00110";
                when x"214D" => data <= "00000";
                when x"214E" => data <= "11001";
                when x"214F" => data <= "00000";
                when x"2150" => data <= "00110";
                when x"2151" => data <= "00110";
                when x"2152" => data <= "00000";
                when x"2153" => data <= "00000";
                when x"2154" => data <= "00110";
                when x"2155" => data <= "00000";
                when x"2156" => data <= "01001";
                when x"2157" => data <= "00000";
                when x"2158" => data <= "00000";
                when x"2159" => data <= "00100";
                when x"215A" => data <= "00110";
                when x"215B" => data <= "00000";
                when x"215C" => data <= "00000";
                when x"215D" => data <= "00110";
                when x"215E" => data <= "00110";
                when x"215F" => data <= "00000";
                when x"2160" => data <= "00000";
                when x"2161" => data <= "11000";
                when x"2162" => data <= "00000";
                when x"2163" => data <= "00000";
                when x"2164" => data <= "00000";
                when x"2165" => data <= "00110";
                when x"2166" => data <= "00110";
                when x"2167" => data <= "00110";
                when x"2168" => data <= "00110";
                when x"2169" => data <= "11011";
                when x"216A" => data <= "00000";
                when x"216B" => data <= "00000";
                when x"216C" => data <= "10110";
                when x"216D" => data <= "00000";
                when x"216E" => data <= "11110";
                when x"216F" => data <= "00110";
                when x"2170" => data <= "00110";
                when x"2171" => data <= "01011";
                when x"2172" => data <= "00000";
                when x"2173" => data <= "00110";
                when x"2174" => data <= "00110";
                when x"2175" => data <= "00110";
                when x"2176" => data <= "00110";
                when x"2177" => data <= "11101";
                when x"2178" => data <= "11001";
                when x"2179" => data <= "00000";
                when x"217A" => data <= "00000";
                when x"217B" => data <= "00110";
                when x"217C" => data <= "00110";
                when x"217D" => data <= "00000";
                when x"217E" => data <= "00110";
                when x"217F" => data <= "00110";
                when x"2180" => data <= "00000";
                when x"2181" => data <= "11000";
                when x"2182" => data <= "01101";
                when x"2183" => data <= "00000";
                when x"2184" => data <= "00000";
                when x"2185" => data <= "00000";
                when x"2186" => data <= "00110";
                when x"2187" => data <= "00110";
                when x"2188" => data <= "00110";
                when x"2189" => data <= "00000";
                when x"218A" => data <= "11001";
                when x"218B" => data <= "00110";
                when x"218C" => data <= "00110";
                when x"218D" => data <= "00110";
                when x"218E" => data <= "00110";
                when x"218F" => data <= "10100";
                when x"2190" => data <= "00000";
                when x"2191" => data <= "00000";
                when x"2192" => data <= "10100";
                when x"2193" => data <= "00000";
                when x"2194" => data <= "00000";
                when x"2195" => data <= "00000";
                when x"2196" => data <= "00110";
                when x"2197" => data <= "01001";
                when x"2198" => data <= "00001";
                when x"2199" => data <= "00000";
                when x"219A" => data <= "00110";
                when x"219B" => data <= "00000";
                when x"219C" => data <= "00110";
                when x"219D" => data <= "00001";
                when x"219E" => data <= "00000";
                when x"219F" => data <= "00000";
                when x"21A0" => data <= "00110";
                when x"21A1" => data <= "00110";
                when x"21A2" => data <= "00010";
                when x"21A3" => data <= "00110";
                when x"21A4" => data <= "00000";
                when x"21A5" => data <= "00110";
                when x"21A6" => data <= "00110";
                when x"21A7" => data <= "00110";
                when x"21A8" => data <= "10111";
                when x"21A9" => data <= "00110";
                when x"21AA" => data <= "00110";
                when x"21AB" => data <= "01011";
                when x"21AC" => data <= "10010";
                when x"21AD" => data <= "00110";
                when x"21AE" => data <= "00000";
                when x"21AF" => data <= "00000";
                when x"21B0" => data <= "00110";
                when x"21B1" => data <= "00110";
                when x"21B2" => data <= "00000";
                when x"21B3" => data <= "00110";
                when x"21B4" => data <= "00000";
                when x"21B5" => data <= "00110";
                when x"21B6" => data <= "01001";
                when x"21B7" => data <= "00110";
                when x"21B8" => data <= "00111";
                when x"21B9" => data <= "00000";
                when x"21BA" => data <= "00110";
                when x"21BB" => data <= "10001";
                when x"21BC" => data <= "00000";
                when x"21BD" => data <= "01011";
                when x"21BE" => data <= "00000";
                when x"21BF" => data <= "00000";
                when x"21C0" => data <= "00110";
                when x"21C1" => data <= "00110";
                when x"21C2" => data <= "00000";
                when x"21C3" => data <= "00110";
                when x"21C4" => data <= "01100";
                when x"21C5" => data <= "00110";
                when x"21C6" => data <= "10001";
                when x"21C7" => data <= "00000";
                when x"21C8" => data <= "00000";
                when x"21C9" => data <= "00110";
                when x"21CA" => data <= "00110";
                when x"21CB" => data <= "11100";
                when x"21CC" => data <= "11010";
                when x"21CD" => data <= "00110";
                when x"21CE" => data <= "00110";
                when x"21CF" => data <= "00000";
                when x"21D0" => data <= "00000";
                when x"21D1" => data <= "00110";
                when x"21D2" => data <= "00110";
                when x"21D3" => data <= "00110";
                when x"21D4" => data <= "00000";
                when x"21D5" => data <= "00000";
                when x"21D6" => data <= "00011";
                when x"21D7" => data <= "00000";
                when x"21D8" => data <= "00110";
                when x"21D9" => data <= "00110";
                when x"21DA" => data <= "00110";
                when x"21DB" => data <= "10001";
                when x"21DC" => data <= "00000";
                when x"21DD" => data <= "00000";
                when x"21DE" => data <= "00110";
                when x"21DF" => data <= "00000";
                when x"21E0" => data <= "00110";
                when x"21E1" => data <= "10010";
                when x"21E2" => data <= "11010";
                when x"21E3" => data <= "00000";
                when x"21E4" => data <= "00000";
                when x"21E5" => data <= "00110";
                when x"21E6" => data <= "00110";
                when x"21E7" => data <= "00110";
                when x"21E8" => data <= "00000";
                when x"21E9" => data <= "00110";
                when x"21EA" => data <= "00110";
                when x"21EB" => data <= "00000";
                when x"21EC" => data <= "00110";
                when x"21ED" => data <= "00110";
                when x"21EE" => data <= "00000";
                when x"21EF" => data <= "00000";
                when x"21F0" => data <= "00000";
                when x"21F1" => data <= "00110";
                when x"21F2" => data <= "00000";
                when x"21F3" => data <= "00110";
                when x"21F4" => data <= "00000";
                when x"21F5" => data <= "00000";
                when x"21F6" => data <= "00000";
                when x"21F7" => data <= "00110";
                when x"21F8" => data <= "00000";
                when x"21F9" => data <= "00000";
                when x"21FA" => data <= "00110";
                when x"21FB" => data <= "00110";
                when x"21FC" => data <= "00000";
                when x"21FD" => data <= "00110";
                when x"21FE" => data <= "01000";
                when x"21FF" => data <= "00000";
                when x"2200" => data <= "00110";
                when x"2201" => data <= "00000";
                when x"2202" => data <= "00110";
                when x"2203" => data <= "00110";
                when x"2204" => data <= "10011";
                when x"2205" => data <= "11000";
                when x"2206" => data <= "00110";
                when x"2207" => data <= "00000";
                when x"2208" => data <= "00000";
                when x"2209" => data <= "00110";
                when x"220A" => data <= "00001";
                when x"220B" => data <= "01101";
                when x"220C" => data <= "00110";
                when x"220D" => data <= "00000";
                when x"220E" => data <= "00000";
                when x"220F" => data <= "11110";
                when x"2210" => data <= "00110";
                when x"2211" => data <= "00110";
                when x"2212" => data <= "11011";
                when x"2213" => data <= "00000";
                when x"2214" => data <= "00110";
                when x"2215" => data <= "00000";
                when x"2216" => data <= "00000";
                when x"2217" => data <= "00000";
                when x"2218" => data <= "00100";
                when x"2219" => data <= "11100";
                when x"221A" => data <= "00000";
                when x"221B" => data <= "00000";
                when x"221C" => data <= "00110";
                when x"221D" => data <= "00110";
                when x"221E" => data <= "00000";
                when x"221F" => data <= "00000";
                when x"2220" => data <= "11111";
                when x"2221" => data <= "00110";
                when x"2222" => data <= "11001";
                when x"2223" => data <= "00110";
                when x"2224" => data <= "11001";
                when x"2225" => data <= "00000";
                when x"2226" => data <= "10010";
                when x"2227" => data <= "00000";
                when x"2228" => data <= "11011";
                when x"2229" => data <= "00000";
                when x"222A" => data <= "00000";
                when x"222B" => data <= "00110";
                when x"222C" => data <= "00110";
                when x"222D" => data <= "00110";
                when x"222E" => data <= "00000";
                when x"222F" => data <= "00000";
                when x"2230" => data <= "11111";
                when x"2231" => data <= "00110";
                when x"2232" => data <= "00110";
                when x"2233" => data <= "00110";
                when x"2234" => data <= "10001";
                when x"2235" => data <= "01101";
                when x"2236" => data <= "00000";
                when x"2237" => data <= "00110";
                when x"2238" => data <= "11010";
                when x"2239" => data <= "00110";
                when x"223A" => data <= "11110";
                when x"223B" => data <= "00000";
                when x"223C" => data <= "00000";
                when x"223D" => data <= "00110";
                when x"223E" => data <= "00110";
                when x"223F" => data <= "00110";
                when x"2240" => data <= "00110";
                when x"2241" => data <= "00000";
                when x"2242" => data <= "00110";
                when x"2243" => data <= "11001";
                when x"2244" => data <= "00000";
                when x"2245" => data <= "00110";
                when x"2246" => data <= "00000";
                when x"2247" => data <= "11001";
                when x"2248" => data <= "00110";
                when x"2249" => data <= "00110";
                when x"224A" => data <= "11111";
                when x"224B" => data <= "11101";
                when x"224C" => data <= "00000";
                when x"224D" => data <= "00000";
                when x"224E" => data <= "00110";
                when x"224F" => data <= "00000";
                when x"2250" => data <= "00000";
                when x"2251" => data <= "00000";
                when x"2252" => data <= "10001";
                when x"2253" => data <= "00000";
                when x"2254" => data <= "00000";
                when x"2255" => data <= "00110";
                when x"2256" => data <= "00110";
                when x"2257" => data <= "00110";
                when x"2258" => data <= "00000";
                when x"2259" => data <= "00110";
                when x"225A" => data <= "00110";
                when x"225B" => data <= "00000";
                when x"225C" => data <= "00110";
                when x"225D" => data <= "00000";
                when x"225E" => data <= "00110";
                when x"225F" => data <= "00000";
                when x"2260" => data <= "01001";
                when x"2261" => data <= "00000";
                when x"2262" => data <= "00000";
                when x"2263" => data <= "00000";
                when x"2264" => data <= "00000";
                when x"2265" => data <= "00000";
                when x"2266" => data <= "00000";
                when x"2267" => data <= "00110";
                when x"2268" => data <= "00000";
                when x"2269" => data <= "00000";
                when x"226A" => data <= "00000";
                when x"226B" => data <= "00110";
                when x"226C" => data <= "10101";
                when x"226D" => data <= "00110";
                when x"226E" => data <= "00000";
                when x"226F" => data <= "00110";
                when x"2270" => data <= "00110";
                when x"2271" => data <= "00000";
                when x"2272" => data <= "00000";
                when x"2273" => data <= "00000";
                when x"2274" => data <= "00000";
                when x"2275" => data <= "01011";
                when x"2276" => data <= "00000";
                when x"2277" => data <= "00110";
                when x"2278" => data <= "00111";
                when x"2279" => data <= "00000";
                when x"227A" => data <= "00000";
                when x"227B" => data <= "00000";
                when x"227C" => data <= "00000";
                when x"227D" => data <= "00110";
                when x"227E" => data <= "11101";
                when x"227F" => data <= "00110";
                when x"2280" => data <= "00000";
                when x"2281" => data <= "00000";
                when x"2282" => data <= "00110";
                when x"2283" => data <= "00110";
                when x"2284" => data <= "00000";
                when x"2285" => data <= "00000";
                when x"2286" => data <= "00000";
                when x"2287" => data <= "10000";
                when x"2288" => data <= "00110";
                when x"2289" => data <= "00110";
                when x"228A" => data <= "00001";
                when x"228B" => data <= "00110";
                when x"228C" => data <= "00110";
                when x"228D" => data <= "11111";
                when x"228E" => data <= "00000";
                when x"228F" => data <= "00000";
                when x"2290" => data <= "00000";
                when x"2291" => data <= "00000";
                when x"2292" => data <= "01000";
                when x"2293" => data <= "00000";
                when x"2294" => data <= "00000";
                when x"2295" => data <= "00000";
                when x"2296" => data <= "00000";
                when x"2297" => data <= "00000";
                when x"2298" => data <= "00110";
                when x"2299" => data <= "00110";
                when x"229A" => data <= "00000";
                when x"229B" => data <= "00000";
                when x"229C" => data <= "00110";
                when x"229D" => data <= "11111";
                when x"229E" => data <= "00000";
                when x"229F" => data <= "01011";
                when x"22A0" => data <= "00000";
                when x"22A1" => data <= "00111";
                when x"22A2" => data <= "00110";
                when x"22A3" => data <= "10010";
                when x"22A4" => data <= "00110";
                when x"22A5" => data <= "00000";
                when x"22A6" => data <= "00110";
                when x"22A7" => data <= "00110";
                when x"22A8" => data <= "00001";
                when x"22A9" => data <= "00110";
                when x"22AA" => data <= "00110";
                when x"22AB" => data <= "00110";
                when x"22AC" => data <= "00000";
                when x"22AD" => data <= "11101";
                when x"22AE" => data <= "00000";
                when x"22AF" => data <= "00110";
                when x"22B0" => data <= "00000";
                when x"22B1" => data <= "11110";
                when x"22B2" => data <= "01010";
                when x"22B3" => data <= "00000";
                when x"22B4" => data <= "00000";
                when x"22B5" => data <= "00000";
                when x"22B6" => data <= "00000";
                when x"22B7" => data <= "00000";
                when x"22B8" => data <= "00110";
                when x"22B9" => data <= "00110";
                when x"22BA" => data <= "00000";
                when x"22BB" => data <= "00110";
                when x"22BC" => data <= "00000";
                when x"22BD" => data <= "00000";
                when x"22BE" => data <= "00111";
                when x"22BF" => data <= "10110";
                when x"22C0" => data <= "00110";
                when x"22C1" => data <= "11100";
                when x"22C2" => data <= "00110";
                when x"22C3" => data <= "00000";
                when x"22C4" => data <= "11100";
                when x"22C5" => data <= "00000";
                when x"22C6" => data <= "11010";
                when x"22C7" => data <= "00000";
                when x"22C8" => data <= "00000";
                when x"22C9" => data <= "10111";
                when x"22CA" => data <= "00110";
                when x"22CB" => data <= "00000";
                when x"22CC" => data <= "00000";
                when x"22CD" => data <= "00000";
                when x"22CE" => data <= "00110";
                when x"22CF" => data <= "00110";
                when x"22D0" => data <= "11010";
                when x"22D1" => data <= "00000";
                when x"22D2" => data <= "00000";
                when x"22D3" => data <= "00110";
                when x"22D4" => data <= "00110";
                when x"22D5" => data <= "00110";
                when x"22D6" => data <= "00000";
                when x"22D7" => data <= "00110";
                when x"22D8" => data <= "00110";
                when x"22D9" => data <= "00110";
                when x"22DA" => data <= "00000";
                when x"22DB" => data <= "00000";
                when x"22DC" => data <= "10000";
                when x"22DD" => data <= "00110";
                when x"22DE" => data <= "00000";
                when x"22DF" => data <= "11000";
                when x"22E0" => data <= "00000";
                when x"22E1" => data <= "00000";
                when x"22E2" => data <= "00110";
                when x"22E3" => data <= "00110";
                when x"22E4" => data <= "00110";
                when x"22E5" => data <= "00000";
                when x"22E6" => data <= "00000";
                when x"22E7" => data <= "01010";
                when x"22E8" => data <= "11001";
                when x"22E9" => data <= "00000";
                when x"22EA" => data <= "00000";
                when x"22EB" => data <= "00000";
                when x"22EC" => data <= "01110";
                when x"22ED" => data <= "00110";
                when x"22EE" => data <= "00100";
                when x"22EF" => data <= "00110";
                when x"22F0" => data <= "00011";
                when x"22F1" => data <= "10100";
                when x"22F2" => data <= "00110";
                when x"22F3" => data <= "11100";
                when x"22F4" => data <= "00000";
                when x"22F5" => data <= "00100";
                when x"22F6" => data <= "00110";
                when x"22F7" => data <= "00000";
                when x"22F8" => data <= "00110";
                when x"22F9" => data <= "00110";
                when x"22FA" => data <= "00110";
                when x"22FB" => data <= "00110";
                when x"22FC" => data <= "11001";
                when x"22FD" => data <= "00110";
                when x"22FE" => data <= "00110";
                when x"22FF" => data <= "00110";
                when x"2300" => data <= "00110";
                when x"2301" => data <= "00110";
                when x"2302" => data <= "00110";
                when x"2303" => data <= "00110";
                when x"2304" => data <= "00101";
                when x"2305" => data <= "10110";
                when x"2306" => data <= "11011";
                when x"2307" => data <= "00110";
                when x"2308" => data <= "00000";
                when x"2309" => data <= "10101";
                when x"230A" => data <= "00000";
                when x"230B" => data <= "00110";
                when x"230C" => data <= "00110";
                when x"230D" => data <= "10010";
                when x"230E" => data <= "00110";
                when x"230F" => data <= "00110";
                when x"2310" => data <= "00110";
                when x"2311" => data <= "00000";
                when x"2312" => data <= "00110";
                when x"2313" => data <= "00000";
                when x"2314" => data <= "00000";
                when x"2315" => data <= "00000";
                when x"2316" => data <= "00000";
                when x"2317" => data <= "01010";
                when x"2318" => data <= "01011";
                when x"2319" => data <= "01101";
                when x"231A" => data <= "00110";
                when x"231B" => data <= "00110";
                when x"231C" => data <= "00110";
                when x"231D" => data <= "00110";
                when x"231E" => data <= "10011";
                when x"231F" => data <= "00000";
                when x"2320" => data <= "00000";
                when x"2321" => data <= "10100";
                when x"2322" => data <= "00110";
                when x"2323" => data <= "00000";
                when x"2324" => data <= "00110";
                when x"2325" => data <= "00110";
                when x"2326" => data <= "10101";
                when x"2327" => data <= "01101";
                when x"2328" => data <= "00110";
                when x"2329" => data <= "00011";
                when x"232A" => data <= "00110";
                when x"232B" => data <= "01111";
                when x"232C" => data <= "00110";
                when x"232D" => data <= "00000";
                when x"232E" => data <= "00000";
                when x"232F" => data <= "00110";
                when x"2330" => data <= "10111";
                when x"2331" => data <= "01111";
                when x"2332" => data <= "00110";
                when x"2333" => data <= "00110";
                when x"2334" => data <= "00000";
                when x"2335" => data <= "00110";
                when x"2336" => data <= "00000";
                when x"2337" => data <= "01110";
                when x"2338" => data <= "00110";
                when x"2339" => data <= "00000";
                when x"233A" => data <= "00110";
                when x"233B" => data <= "00110";
                when x"233C" => data <= "00000";
                when x"233D" => data <= "00111";
                when x"233E" => data <= "00110";
                when x"233F" => data <= "11011";
                when x"2340" => data <= "01101";
                when x"2341" => data <= "01011";
                when x"2342" => data <= "00110";
                when x"2343" => data <= "11010";
                when x"2344" => data <= "00110";
                when x"2345" => data <= "00000";
                when x"2346" => data <= "00000";
                when x"2347" => data <= "00110";
                when x"2348" => data <= "01101";
                when x"2349" => data <= "00110";
                when x"234A" => data <= "00000";
                when x"234B" => data <= "00110";
                when x"234C" => data <= "00110";
                when x"234D" => data <= "00110";
                when x"234E" => data <= "00000";
                when x"234F" => data <= "00110";
                when x"2350" => data <= "11101";
                when x"2351" => data <= "00110";
                when x"2352" => data <= "01001";
                when x"2353" => data <= "00000";
                when x"2354" => data <= "00000";
                when x"2355" => data <= "00000";
                when x"2356" => data <= "00000";
                when x"2357" => data <= "00110";
                when x"2358" => data <= "00110";
                when x"2359" => data <= "00110";
                when x"235A" => data <= "00110";
                when x"235B" => data <= "11001";
                when x"235C" => data <= "00110";
                when x"235D" => data <= "00110";
                when x"235E" => data <= "00000";
                when x"235F" => data <= "00110";
                when x"2360" => data <= "00110";
                when x"2361" => data <= "00110";
                when x"2362" => data <= "00110";
                when x"2363" => data <= "00110";
                when x"2364" => data <= "00000";
                when x"2365" => data <= "00000";
                when x"2366" => data <= "00000";
                when x"2367" => data <= "00110";
                when x"2368" => data <= "00000";
                when x"2369" => data <= "10011";
                when x"236A" => data <= "00000";
                when x"236B" => data <= "00000";
                when x"236C" => data <= "11110";
                when x"236D" => data <= "00110";
                when x"236E" => data <= "00000";
                when x"236F" => data <= "11010";
                when x"2370" => data <= "00110";
                when x"2371" => data <= "01010";
                when x"2372" => data <= "10101";
                when x"2373" => data <= "01110";
                when x"2374" => data <= "00000";
                when x"2375" => data <= "00001";
                when x"2376" => data <= "00000";
                when x"2377" => data <= "00000";
                when x"2378" => data <= "00000";
                when x"2379" => data <= "00110";
                when x"237A" => data <= "00000";
                when x"237B" => data <= "01011";
                when x"237C" => data <= "00110";
                when x"237D" => data <= "00000";
                when x"237E" => data <= "00110";
                when x"237F" => data <= "00000";
                when x"2380" => data <= "00110";
                when x"2381" => data <= "00110";
                when x"2382" => data <= "00000";
                when x"2383" => data <= "01101";
                when x"2384" => data <= "00110";
                when x"2385" => data <= "11001";
                when x"2386" => data <= "00110";
                when x"2387" => data <= "00000";
                when x"2388" => data <= "00110";
                when x"2389" => data <= "00000";
                when x"238A" => data <= "00110";
                when x"238B" => data <= "00110";
                when x"238C" => data <= "00110";
                when x"238D" => data <= "00000";
                when x"238E" => data <= "00000";
                when x"238F" => data <= "00000";
                when x"2390" => data <= "00110";
                when x"2391" => data <= "00110";
                when x"2392" => data <= "00110";
                when x"2393" => data <= "00000";
                when x"2394" => data <= "00000";
                when x"2395" => data <= "00000";
                when x"2396" => data <= "00110";
                when x"2397" => data <= "11111";
                when x"2398" => data <= "11000";
                when x"2399" => data <= "00110";
                when x"239A" => data <= "00000";
                when x"239B" => data <= "10101";
                when x"239C" => data <= "00000";
                when x"239D" => data <= "01100";
                when x"239E" => data <= "00000";
                when x"239F" => data <= "00000";
                when x"23A0" => data <= "00110";
                when x"23A1" => data <= "00000";
                when x"23A2" => data <= "00110";
                when x"23A3" => data <= "00000";
                when x"23A4" => data <= "00000";
                when x"23A5" => data <= "00110";
                when x"23A6" => data <= "00000";
                when x"23A7" => data <= "00110";
                when x"23A8" => data <= "01001";
                when x"23A9" => data <= "00110";
                when x"23AA" => data <= "00110";
                when x"23AB" => data <= "00000";
                when x"23AC" => data <= "00110";
                when x"23AD" => data <= "00010";
                when x"23AE" => data <= "00110";
                when x"23AF" => data <= "00110";
                when x"23B0" => data <= "00110";
                when x"23B1" => data <= "01011";
                when x"23B2" => data <= "00000";
                when x"23B3" => data <= "00110";
                when x"23B4" => data <= "00000";
                when x"23B5" => data <= "01100";
                when x"23B6" => data <= "00000";
                when x"23B7" => data <= "00000";
                when x"23B8" => data <= "10011";
                when x"23B9" => data <= "00110";
                when x"23BA" => data <= "00110";
                when x"23BB" => data <= "00011";
                when x"23BC" => data <= "00000";
                when x"23BD" => data <= "00110";
                when x"23BE" => data <= "00110";
                when x"23BF" => data <= "00110";
                when x"23C0" => data <= "00110";
                when x"23C1" => data <= "00110";
                when x"23C2" => data <= "00110";
                when x"23C3" => data <= "00000";
                when x"23C4" => data <= "00110";
                when x"23C5" => data <= "00000";
                when x"23C6" => data <= "01000";
                when x"23C7" => data <= "10011";
                when x"23C8" => data <= "00110";
                when x"23C9" => data <= "00110";
                when x"23CA" => data <= "00000";
                when x"23CB" => data <= "00110";
                when x"23CC" => data <= "00000";
                when x"23CD" => data <= "00110";
                when x"23CE" => data <= "00000";
                when x"23CF" => data <= "00110";
                when x"23D0" => data <= "00000";
                when x"23D1" => data <= "00110";
                when x"23D2" => data <= "00000";
                when x"23D3" => data <= "11111";
                when x"23D4" => data <= "11100";
                when x"23D5" => data <= "00110";
                when x"23D6" => data <= "00110";
                when x"23D7" => data <= "00000";
                when x"23D8" => data <= "00000";
                when x"23D9" => data <= "01101";
                when x"23DA" => data <= "00000";
                when x"23DB" => data <= "10101";
                when x"23DC" => data <= "00000";
                when x"23DD" => data <= "00000";
                when x"23DE" => data <= "00000";
                when x"23DF" => data <= "00110";
                when x"23E0" => data <= "00000";
                when x"23E1" => data <= "00110";
                when x"23E2" => data <= "00110";
                when x"23E3" => data <= "00110";
                when x"23E4" => data <= "00000";
                when x"23E5" => data <= "01111";
                when x"23E6" => data <= "00110";
                when x"23E7" => data <= "01011";
                when x"23E8" => data <= "00110";
                when x"23E9" => data <= "00000";
                when x"23EA" => data <= "00000";
                when x"23EB" => data <= "00110";
                when x"23EC" => data <= "00000";
                when x"23ED" => data <= "00000";
                when x"23EE" => data <= "00000";
                when x"23EF" => data <= "00000";
                when x"23F0" => data <= "11010";
                when x"23F1" => data <= "00000";
                when x"23F2" => data <= "00110";
                when x"23F3" => data <= "00110";
                when x"23F4" => data <= "00000";
                when x"23F5" => data <= "00000";
                when x"23F6" => data <= "00000";
                when x"23F7" => data <= "00000";
                when x"23F8" => data <= "00000";
                when x"23F9" => data <= "00110";
                when x"23FA" => data <= "00110";
                when x"23FB" => data <= "01011";
                when x"23FC" => data <= "00000";
                when x"23FD" => data <= "00000";
                when x"23FE" => data <= "01011";
                when x"23FF" => data <= "00110";
                when x"2400" => data <= "00110";
                when x"2401" => data <= "00000";
                when x"2402" => data <= "00000";
                when x"2403" => data <= "00000";
                when x"2404" => data <= "00110";
                when x"2405" => data <= "00000";
                when x"2406" => data <= "00000";
                when x"2407" => data <= "00000";
                when x"2408" => data <= "00110";
                when x"2409" => data <= "00110";
                when x"240A" => data <= "10111";
                when x"240B" => data <= "00110";
                when x"240C" => data <= "00110";
                when x"240D" => data <= "10101";
                when x"240E" => data <= "10000";
                when x"240F" => data <= "00000";
                when x"2410" => data <= "01001";
                when x"2411" => data <= "01000";
                when x"2412" => data <= "00000";
                when x"2413" => data <= "00000";
                when x"2414" => data <= "00000";
                when x"2415" => data <= "00110";
                when x"2416" => data <= "00000";
                when x"2417" => data <= "00110";
                when x"2418" => data <= "00101";
                when x"2419" => data <= "01101";
                when x"241A" => data <= "00110";
                when x"241B" => data <= "01011";
                when x"241C" => data <= "00000";
                when x"241D" => data <= "10010";
                when x"241E" => data <= "10000";
                when x"241F" => data <= "00110";
                when x"2420" => data <= "11111";
                when x"2421" => data <= "00000";
                when x"2422" => data <= "00110";
                when x"2423" => data <= "00110";
                when x"2424" => data <= "00000";
                when x"2425" => data <= "00000";
                when x"2426" => data <= "00110";
                when x"2427" => data <= "00000";
                when x"2428" => data <= "00110";
                when x"2429" => data <= "00110";
                when x"242A" => data <= "00001";
                when x"242B" => data <= "00110";
                when x"242C" => data <= "00110";
                when x"242D" => data <= "00110";
                when x"242E" => data <= "00110";
                when x"242F" => data <= "00000";
                when x"2430" => data <= "10101";
                when x"2431" => data <= "00110";
                when x"2432" => data <= "00000";
                when x"2433" => data <= "00000";
                when x"2434" => data <= "00110";
                when x"2435" => data <= "00000";
                when x"2436" => data <= "01010";
                when x"2437" => data <= "00000";
                when x"2438" => data <= "00110";
                when x"2439" => data <= "00000";
                when x"243A" => data <= "00000";
                when x"243B" => data <= "00110";
                when x"243C" => data <= "00000";
                when x"243D" => data <= "00000";
                when x"243E" => data <= "00000";
                when x"243F" => data <= "00000";
                when x"2440" => data <= "00110";
                when x"2441" => data <= "00000";
                when x"2442" => data <= "00000";
                when x"2443" => data <= "00110";
                when x"2444" => data <= "00000";
                when x"2445" => data <= "00110";
                when x"2446" => data <= "00000";
                when x"2447" => data <= "00000";
                when x"2448" => data <= "00110";
                when x"2449" => data <= "00000";
                when x"244A" => data <= "00110";
                when x"244B" => data <= "00110";
                when x"244C" => data <= "00000";
                when x"244D" => data <= "00000";
                when x"244E" => data <= "00110";
                when x"244F" => data <= "00110";
                when x"2450" => data <= "01111";
                when x"2451" => data <= "00110";
                when x"2452" => data <= "00000";
                when x"2453" => data <= "01100";
                when x"2454" => data <= "01101";
                when x"2455" => data <= "10101";
                when x"2456" => data <= "00000";
                when x"2457" => data <= "00110";
                when x"2458" => data <= "00110";
                when x"2459" => data <= "10000";
                when x"245A" => data <= "00010";
                when x"245B" => data <= "00000";
                when x"245C" => data <= "10010";
                when x"245D" => data <= "00000";
                when x"245E" => data <= "00110";
                when x"245F" => data <= "01110";
                when x"2460" => data <= "00111";
                when x"2461" => data <= "00110";
                when x"2462" => data <= "00110";
                when x"2463" => data <= "00000";
                when x"2464" => data <= "00000";
                when x"2465" => data <= "10110";
                when x"2466" => data <= "00000";
                when x"2467" => data <= "00000";
                when x"2468" => data <= "00110";
                when x"2469" => data <= "00110";
                when x"246A" => data <= "00110";
                when x"246B" => data <= "00000";
                when x"246C" => data <= "00000";
                when x"246D" => data <= "00000";
                when x"246E" => data <= "10101";
                when x"246F" => data <= "00000";
                when x"2470" => data <= "00000";
                when x"2471" => data <= "10101";
                when x"2472" => data <= "00000";
                when x"2473" => data <= "00000";
                when x"2474" => data <= "10111";
                when x"2475" => data <= "00000";
                when x"2476" => data <= "00110";
                when x"2477" => data <= "00000";
                when x"2478" => data <= "00110";
                when x"2479" => data <= "00000";
                when x"247A" => data <= "00000";
                when x"247B" => data <= "00000";
                when x"247C" => data <= "00110";
                when x"247D" => data <= "00000";
                when x"247E" => data <= "01101";
                when x"247F" => data <= "00110";
                when x"2480" => data <= "11100";
                when x"2481" => data <= "00110";
                when x"2482" => data <= "00110";
                when x"2483" => data <= "00000";
                when x"2484" => data <= "00000";
                when x"2485" => data <= "00000";
                when x"2486" => data <= "00000";
                when x"2487" => data <= "00000";
                when x"2488" => data <= "00000";
                when x"2489" => data <= "01001";
                when x"248A" => data <= "00000";
                when x"248B" => data <= "00000";
                when x"248C" => data <= "00000";
                when x"248D" => data <= "00110";
                when x"248E" => data <= "00110";
                when x"248F" => data <= "01010";
                when x"2490" => data <= "00000";
                when x"2491" => data <= "00000";
                when x"2492" => data <= "00110";
                when x"2493" => data <= "00110";
                when x"2494" => data <= "00110";
                when x"2495" => data <= "00110";
                when x"2496" => data <= "00110";
                when x"2497" => data <= "00000";
                when x"2498" => data <= "00110";
                when x"2499" => data <= "00000";
                when x"249A" => data <= "00000";
                when x"249B" => data <= "00110";
                when x"249C" => data <= "00110";
                when x"249D" => data <= "00110";
                when x"249E" => data <= "00000";
                when x"249F" => data <= "00000";
                when x"24A0" => data <= "00110";
                when x"24A1" => data <= "00110";
                when x"24A2" => data <= "10111";
                when x"24A3" => data <= "00000";
                when x"24A4" => data <= "11000";
                when x"24A5" => data <= "00110";
                when x"24A6" => data <= "00000";
                when x"24A7" => data <= "00000";
                when x"24A8" => data <= "00110";
                when x"24A9" => data <= "00110";
                when x"24AA" => data <= "00110";
                when x"24AB" => data <= "00000";
                when x"24AC" => data <= "00000";
                when x"24AD" => data <= "01010";
                when x"24AE" => data <= "01011";
                when x"24AF" => data <= "00000";
                when x"24B0" => data <= "00110";
                when x"24B1" => data <= "00110";
                when x"24B2" => data <= "10110";
                when x"24B3" => data <= "10111";
                when x"24B4" => data <= "10010";
                when x"24B5" => data <= "00110";
                when x"24B6" => data <= "00110";
                when x"24B7" => data <= "11010";
                when x"24B8" => data <= "00110";
                when x"24B9" => data <= "00000";
                when x"24BA" => data <= "00000";
                when x"24BB" => data <= "00000";
                when x"24BC" => data <= "11110";
                when x"24BD" => data <= "00000";
                when x"24BE" => data <= "00000";
                when x"24BF" => data <= "00000";
                when x"24C0" => data <= "10010";
                when x"24C1" => data <= "00000";
                when x"24C2" => data <= "00000";
                when x"24C3" => data <= "00000";
                when x"24C4" => data <= "00000";
                when x"24C5" => data <= "00110";
                when x"24C6" => data <= "00110";
                when x"24C7" => data <= "00000";
                when x"24C8" => data <= "00000";
                when x"24C9" => data <= "00000";
                when x"24CA" => data <= "01010";
                when x"24CB" => data <= "00000";
                when x"24CC" => data <= "11001";
                when x"24CD" => data <= "00110";
                when x"24CE" => data <= "00110";
                when x"24CF" => data <= "00110";
                when x"24D0" => data <= "00000";
                when x"24D1" => data <= "00000";
                when x"24D2" => data <= "01111";
                when x"24D3" => data <= "00010";
                when x"24D4" => data <= "00110";
                when x"24D5" => data <= "00000";
                when x"24D6" => data <= "10001";
                when x"24D7" => data <= "00000";
                when x"24D8" => data <= "00000";
                when x"24D9" => data <= "00000";
                when x"24DA" => data <= "00110";
                when x"24DB" => data <= "00000";
                when x"24DC" => data <= "00110";
                when x"24DD" => data <= "00110";
                when x"24DE" => data <= "00000";
                when x"24DF" => data <= "00110";
                when x"24E0" => data <= "00110";
                when x"24E1" => data <= "00000";
                when x"24E2" => data <= "01011";
                when x"24E3" => data <= "10111";
                when x"24E4" => data <= "11100";
                when x"24E5" => data <= "00000";
                when x"24E6" => data <= "01100";
                when x"24E7" => data <= "11001";
                when x"24E8" => data <= "00000";
                when x"24E9" => data <= "00110";
                when x"24EA" => data <= "00110";
                when x"24EB" => data <= "00000";
                when x"24EC" => data <= "00000";
                when x"24ED" => data <= "00110";
                when x"24EE" => data <= "01101";
                when x"24EF" => data <= "00110";
                when x"24F0" => data <= "00000";
                when x"24F1" => data <= "10101";
                when x"24F2" => data <= "00000";
                when x"24F3" => data <= "00110";
                when x"24F4" => data <= "00000";
                when x"24F5" => data <= "00110";
                when x"24F6" => data <= "00000";
                when x"24F7" => data <= "00110";
                when x"24F8" => data <= "00110";
                when x"24F9" => data <= "00110";
                when x"24FA" => data <= "00000";
                when x"24FB" => data <= "00110";
                when x"24FC" => data <= "01111";
                when x"24FD" => data <= "00110";
                when x"24FE" => data <= "00000";
                when x"24FF" => data <= "11100";
                when x"2500" => data <= "11000";
                when x"2501" => data <= "00110";
                when x"2502" => data <= "00110";
                when x"2503" => data <= "00110";
                when x"2504" => data <= "01101";
                when x"2505" => data <= "11100";
                when x"2506" => data <= "00000";
                when x"2507" => data <= "00110";
                when x"2508" => data <= "00101";
                when x"2509" => data <= "01111";
                when x"250A" => data <= "00110";
                when x"250B" => data <= "00000";
                when x"250C" => data <= "00110";
                when x"250D" => data <= "00000";
                when x"250E" => data <= "00000";
                when x"250F" => data <= "00000";
                when x"2510" => data <= "00110";
                when x"2511" => data <= "00000";
                when x"2512" => data <= "00000";
                when x"2513" => data <= "10011";
                when x"2514" => data <= "00110";
                when x"2515" => data <= "11000";
                when x"2516" => data <= "00000";
                when x"2517" => data <= "00000";
                when x"2518" => data <= "00000";
                when x"2519" => data <= "00110";
                when x"251A" => data <= "01110";
                when x"251B" => data <= "00110";
                when x"251C" => data <= "00000";
                when x"251D" => data <= "01001";
                when x"251E" => data <= "00000";
                when x"251F" => data <= "00000";
                when x"2520" => data <= "01110";
                when x"2521" => data <= "00110";
                when x"2522" => data <= "01000";
                when x"2523" => data <= "01110";
                when x"2524" => data <= "00110";
                when x"2525" => data <= "00000";
                when x"2526" => data <= "00000";
                when x"2527" => data <= "00000";
                when x"2528" => data <= "00000";
                when x"2529" => data <= "00000";
                when x"252A" => data <= "00110";
                when x"252B" => data <= "11000";
                when x"252C" => data <= "00000";
                when x"252D" => data <= "00110";
                when x"252E" => data <= "00111";
                when x"252F" => data <= "00110";
                when x"2530" => data <= "00000";
                when x"2531" => data <= "00000";
                when x"2532" => data <= "11100";
                when x"2533" => data <= "00110";
                when x"2534" => data <= "00000";
                when x"2535" => data <= "10001";
                when x"2536" => data <= "00110";
                when x"2537" => data <= "10110";
                when x"2538" => data <= "00000";
                when x"2539" => data <= "00000";
                when x"253A" => data <= "00110";
                when x"253B" => data <= "00110";
                when x"253C" => data <= "01110";
                when x"253D" => data <= "00000";
                when x"253E" => data <= "00110";
                when x"253F" => data <= "00110";
                when x"2540" => data <= "00000";
                when x"2541" => data <= "00110";
                when x"2542" => data <= "11100";
                when x"2543" => data <= "10011";
                when x"2544" => data <= "11111";
                when x"2545" => data <= "01111";
                when x"2546" => data <= "00000";
                when x"2547" => data <= "00110";
                when x"2548" => data <= "00000";
                when x"2549" => data <= "00110";
                when x"254A" => data <= "00110";
                when x"254B" => data <= "00110";
                when x"254C" => data <= "01111";
                when x"254D" => data <= "00110";
                when x"254E" => data <= "00000";
                when x"254F" => data <= "00000";
                when x"2550" => data <= "00110";
                when x"2551" => data <= "00110";
                when x"2552" => data <= "00110";
                when x"2553" => data <= "00000";
                when x"2554" => data <= "00110";
                when x"2555" => data <= "00110";
                when x"2556" => data <= "00000";
                when x"2557" => data <= "01101";
                when x"2558" => data <= "00000";
                when x"2559" => data <= "00110";
                when x"255A" => data <= "00110";
                when x"255B" => data <= "00000";
                when x"255C" => data <= "00110";
                when x"255D" => data <= "00000";
                when x"255E" => data <= "00110";
                when x"255F" => data <= "00000";
                when x"2560" => data <= "00110";
                when x"2561" => data <= "00110";
                when x"2562" => data <= "00000";
                when x"2563" => data <= "00110";
                when x"2564" => data <= "00110";
                when x"2565" => data <= "01101";
                when x"2566" => data <= "10101";
                when x"2567" => data <= "00000";
                when x"2568" => data <= "10000";
                when x"2569" => data <= "00110";
                when x"256A" => data <= "00000";
                when x"256B" => data <= "00000";
                when x"256C" => data <= "00110";
                when x"256D" => data <= "00110";
                when x"256E" => data <= "00110";
                when x"256F" => data <= "00000";
                when x"2570" => data <= "10011";
                when x"2571" => data <= "00000";
                when x"2572" => data <= "00110";
                when x"2573" => data <= "00000";
                when x"2574" => data <= "01011";
                when x"2575" => data <= "00110";
                when x"2576" => data <= "00110";
                when x"2577" => data <= "00000";
                when x"2578" => data <= "00110";
                when x"2579" => data <= "00000";
                when x"257A" => data <= "00000";
                when x"257B" => data <= "00000";
                when x"257C" => data <= "01101";
                when x"257D" => data <= "11100";
                when x"257E" => data <= "11110";
                when x"257F" => data <= "00110";
                when x"2580" => data <= "00000";
                when x"2581" => data <= "00110";
                when x"2582" => data <= "00000";
                when x"2583" => data <= "00000";
                when x"2584" => data <= "00000";
                when x"2585" => data <= "00001";
                when x"2586" => data <= "00110";
                when x"2587" => data <= "00000";
                when x"2588" => data <= "00110";
                when x"2589" => data <= "00000";
                when x"258A" => data <= "00110";
                when x"258B" => data <= "00110";
                when x"258C" => data <= "01101";
                when x"258D" => data <= "00110";
                when x"258E" => data <= "11000";
                when x"258F" => data <= "00110";
                when x"2590" => data <= "00000";
                when x"2591" => data <= "00110";
                when x"2592" => data <= "00110";
                when x"2593" => data <= "00110";
                when x"2594" => data <= "00110";
                when x"2595" => data <= "01111";
                when x"2596" => data <= "00110";
                when x"2597" => data <= "00110";
                when x"2598" => data <= "00000";
                when x"2599" => data <= "10111";
                when x"259A" => data <= "00110";
                when x"259B" => data <= "00110";
                when x"259C" => data <= "00110";
                when x"259D" => data <= "11111";
                when x"259E" => data <= "00110";
                when x"259F" => data <= "00000";
                when x"25A0" => data <= "00000";
                when x"25A1" => data <= "11100";
                when x"25A2" => data <= "00110";
                when x"25A3" => data <= "00000";
                when x"25A4" => data <= "00000";
                when x"25A5" => data <= "00110";
                when x"25A6" => data <= "00110";
                when x"25A7" => data <= "11000";
                when x"25A8" => data <= "00000";
                when x"25A9" => data <= "00110";
                when x"25AA" => data <= "00110";
                when x"25AB" => data <= "10101";
                when x"25AC" => data <= "00000";
                when x"25AD" => data <= "11001";
                when x"25AE" => data <= "00110";
                when x"25AF" => data <= "00000";
                when x"25B0" => data <= "00110";
                when x"25B1" => data <= "00110";
                when x"25B2" => data <= "00000";
                when x"25B3" => data <= "00110";
                when x"25B4" => data <= "10100";
                when x"25B5" => data <= "00000";
                when x"25B6" => data <= "01100";
                when x"25B7" => data <= "00110";
                when x"25B8" => data <= "11010";
                when x"25B9" => data <= "00000";
                when x"25BA" => data <= "00110";
                when x"25BB" => data <= "00110";
                when x"25BC" => data <= "00110";
                when x"25BD" => data <= "00110";
                when x"25BE" => data <= "00110";
                when x"25BF" => data <= "00000";
                when x"25C0" => data <= "00110";
                when x"25C1" => data <= "11100";
                when x"25C2" => data <= "00110";
                when x"25C3" => data <= "00000";
                when x"25C4" => data <= "00011";
                when x"25C5" => data <= "11100";
                when x"25C6" => data <= "11110";
                when x"25C7" => data <= "01101";
                when x"25C8" => data <= "00000";
                when x"25C9" => data <= "00000";
                when x"25CA" => data <= "11111";
                when x"25CB" => data <= "00000";
                when x"25CC" => data <= "00110";
                when x"25CD" => data <= "00110";
                when x"25CE" => data <= "10111";
                when x"25CF" => data <= "00000";
                when x"25D0" => data <= "00110";
                when x"25D1" => data <= "00000";
                when x"25D2" => data <= "00000";
                when x"25D3" => data <= "00110";
                when x"25D4" => data <= "00110";
                when x"25D5" => data <= "00000";
                when x"25D6" => data <= "00000";
                when x"25D7" => data <= "11001";
                when x"25D8" => data <= "00000";
                when x"25D9" => data <= "01100";
                when x"25DA" => data <= "00110";
                when x"25DB" => data <= "00000";
                when x"25DC" => data <= "00110";
                when x"25DD" => data <= "00000";
                when x"25DE" => data <= "00111";
                when x"25DF" => data <= "00110";
                when x"25E0" => data <= "00000";
                when x"25E1" => data <= "00110";
                when x"25E2" => data <= "00000";
                when x"25E3" => data <= "11000";
                when x"25E4" => data <= "00110";
                when x"25E5" => data <= "00000";
                when x"25E6" => data <= "10100";
                when x"25E7" => data <= "00000";
                when x"25E8" => data <= "00110";
                when x"25E9" => data <= "00110";
                when x"25EA" => data <= "00110";
                when x"25EB" => data <= "00110";
                when x"25EC" => data <= "11101";
                when x"25ED" => data <= "00000";
                when x"25EE" => data <= "00000";
                when x"25EF" => data <= "00000";
                when x"25F0" => data <= "00110";
                when x"25F1" => data <= "00000";
                when x"25F2" => data <= "00000";
                when x"25F3" => data <= "01110";
                when x"25F4" => data <= "00000";
                when x"25F5" => data <= "00110";
                when x"25F6" => data <= "00000";
                when x"25F7" => data <= "00000";
                when x"25F8" => data <= "00110";
                when x"25F9" => data <= "00110";
                when x"25FA" => data <= "00000";
                when x"25FB" => data <= "00110";
                when x"25FC" => data <= "00110";
                when x"25FD" => data <= "00111";
                when x"25FE" => data <= "01101";
                when x"25FF" => data <= "00000";
                when x"2600" => data <= "00000";
                when x"2601" => data <= "00110";
                when x"2602" => data <= "00110";
                when x"2603" => data <= "00110";
                when x"2604" => data <= "00110";
                when x"2605" => data <= "01101";
                when x"2606" => data <= "00110";
                when x"2607" => data <= "00001";
                when x"2608" => data <= "00110";
                when x"2609" => data <= "00110";
                when x"260A" => data <= "00110";
                when x"260B" => data <= "00001";
                when x"260C" => data <= "00000";
                when x"260D" => data <= "00110";
                when x"260E" => data <= "00000";
                when x"260F" => data <= "00110";
                when x"2610" => data <= "10101";
                when x"2611" => data <= "00000";
                when x"2612" => data <= "00000";
                when x"2613" => data <= "11110";
                when x"2614" => data <= "00011";
                when x"2615" => data <= "00110";
                when x"2616" => data <= "01001";
                when x"2617" => data <= "01001";
                when x"2618" => data <= "00110";
                when x"2619" => data <= "00110";
                when x"261A" => data <= "00110";
                when x"261B" => data <= "00000";
                when x"261C" => data <= "00010";
                when x"261D" => data <= "01110";
                when x"261E" => data <= "00110";
                when x"261F" => data <= "00000";
                when x"2620" => data <= "00110";
                when x"2621" => data <= "00110";
                when x"2622" => data <= "00000";
                when x"2623" => data <= "11100";
                when x"2624" => data <= "00110";
                when x"2625" => data <= "00110";
                when x"2626" => data <= "00000";
                when x"2627" => data <= "00000";
                when x"2628" => data <= "00110";
                when x"2629" => data <= "00000";
                when x"262A" => data <= "00110";
                when x"262B" => data <= "00101";
                when x"262C" => data <= "00110";
                when x"262D" => data <= "00000";
                when x"262E" => data <= "00000";
                when x"262F" => data <= "10111";
                when x"2630" => data <= "00110";
                when x"2631" => data <= "11011";
                when x"2632" => data <= "11100";
                when x"2633" => data <= "01110";
                when x"2634" => data <= "00000";
                when x"2635" => data <= "00000";
                when x"2636" => data <= "00110";
                when x"2637" => data <= "00000";
                when x"2638" => data <= "00000";
                when x"2639" => data <= "00110";
                when x"263A" => data <= "00000";
                when x"263B" => data <= "00000";
                when x"263C" => data <= "00110";
                when x"263D" => data <= "00110";
                when x"263E" => data <= "11111";
                when x"263F" => data <= "00101";
                when x"2640" => data <= "00110";
                when x"2641" => data <= "01101";
                when x"2642" => data <= "01011";
                when x"2643" => data <= "00110";
                when x"2644" => data <= "01110";
                when x"2645" => data <= "00000";
                when x"2646" => data <= "00110";
                when x"2647" => data <= "00000";
                when x"2648" => data <= "00110";
                when x"2649" => data <= "00110";
                when x"264A" => data <= "00110";
                when x"264B" => data <= "00110";
                when x"264C" => data <= "00110";
                when x"264D" => data <= "00000";
                when x"264E" => data <= "00110";
                when x"264F" => data <= "11111";
                when x"2650" => data <= "00110";
                when x"2651" => data <= "00000";
                when x"2652" => data <= "00000";
                when x"2653" => data <= "00000";
                when x"2654" => data <= "00110";
                when x"2655" => data <= "00000";
                when x"2656" => data <= "00000";
                when x"2657" => data <= "00110";
                when x"2658" => data <= "00110";
                when x"2659" => data <= "00110";
                when x"265A" => data <= "00000";
                when x"265B" => data <= "00110";
                when x"265C" => data <= "00110";
                when x"265D" => data <= "00000";
                when x"265E" => data <= "00110";
                when x"265F" => data <= "01010";
                when x"2660" => data <= "00000";
                when x"2661" => data <= "00000";
                when x"2662" => data <= "01101";
                when x"2663" => data <= "11110";
                when x"2664" => data <= "00000";
                when x"2665" => data <= "00000";
                when x"2666" => data <= "01101";
                when x"2667" => data <= "10110";
                when x"2668" => data <= "00000";
                when x"2669" => data <= "00110";
                when x"266A" => data <= "00110";
                when x"266B" => data <= "00000";
                when x"266C" => data <= "10110";
                when x"266D" => data <= "01111";
                when x"266E" => data <= "00000";
                when x"266F" => data <= "00000";
                when x"2670" => data <= "10011";
                when x"2671" => data <= "00100";
                when x"2672" => data <= "00000";
                when x"2673" => data <= "00110";
                when x"2674" => data <= "11000";
                when x"2675" => data <= "00110";
                when x"2676" => data <= "11010";
                when x"2677" => data <= "00000";
                when x"2678" => data <= "00110";
                when x"2679" => data <= "00111";
                when x"267A" => data <= "00110";
                when x"267B" => data <= "00000";
                when x"267C" => data <= "00110";
                when x"267D" => data <= "10011";
                when x"267E" => data <= "00110";
                when x"267F" => data <= "00110";
                when x"2680" => data <= "01011";
                when x"2681" => data <= "00000";
                when x"2682" => data <= "00110";
                when x"2683" => data <= "01111";
                when x"2684" => data <= "00101";
                when x"2685" => data <= "00000";
                when x"2686" => data <= "00110";
                when x"2687" => data <= "00000";
                when x"2688" => data <= "00110";
                when x"2689" => data <= "01011";
                when x"268A" => data <= "00110";
                when x"268B" => data <= "00110";
                when x"268C" => data <= "01111";
                when x"268D" => data <= "00110";
                when x"268E" => data <= "00110";
                when x"268F" => data <= "00000";
                when x"2690" => data <= "00001";
                when x"2691" => data <= "01000";
                when x"2692" => data <= "00110";
                when x"2693" => data <= "00000";
                when x"2694" => data <= "00110";
                when x"2695" => data <= "01011";
                when x"2696" => data <= "01000";
                when x"2697" => data <= "00110";
                when x"2698" => data <= "00000";
                when x"2699" => data <= "00000";
                when x"269A" => data <= "00000";
                when x"269B" => data <= "00110";
                when x"269C" => data <= "00000";
                when x"269D" => data <= "00000";
                when x"269E" => data <= "00110";
                when x"269F" => data <= "00000";
                when x"26A0" => data <= "00000";
                when x"26A1" => data <= "00001";
                when x"26A2" => data <= "00110";
                when x"26A3" => data <= "11111";
                when x"26A4" => data <= "00111";
                when x"26A5" => data <= "00000";
                when x"26A6" => data <= "11000";
                when x"26A7" => data <= "00110";
                when x"26A8" => data <= "01101";
                when x"26A9" => data <= "00000";
                when x"26AA" => data <= "00110";
                when x"26AB" => data <= "00000";
                when x"26AC" => data <= "00000";
                when x"26AD" => data <= "00110";
                when x"26AE" => data <= "00000";
                when x"26AF" => data <= "11010";
                when x"26B0" => data <= "00000";
                when x"26B1" => data <= "00110";
                when x"26B2" => data <= "00100";
                when x"26B3" => data <= "11000";
                when x"26B4" => data <= "00000";
                when x"26B5" => data <= "00000";
                when x"26B6" => data <= "10111";
                when x"26B7" => data <= "00000";
                when x"26B8" => data <= "00110";
                when x"26B9" => data <= "00000";
                when x"26BA" => data <= "00000";
                when x"26BB" => data <= "00110";
                when x"26BC" => data <= "10010";
                when x"26BD" => data <= "00110";
                when x"26BE" => data <= "00110";
                when x"26BF" => data <= "00110";
                when x"26C0" => data <= "00000";
                when x"26C1" => data <= "00110";
                when x"26C2" => data <= "01101";
                when x"26C3" => data <= "00000";
                when x"26C4" => data <= "10101";
                when x"26C5" => data <= "00000";
                when x"26C6" => data <= "00000";
                when x"26C7" => data <= "00110";
                when x"26C8" => data <= "11010";
                when x"26C9" => data <= "00110";
                when x"26CA" => data <= "00101";
                when x"26CB" => data <= "00110";
                when x"26CC" => data <= "00000";
                when x"26CD" => data <= "11111";
                when x"26CE" => data <= "01101";
                when x"26CF" => data <= "00000";
                when x"26D0" => data <= "00110";
                when x"26D1" => data <= "00000";
                when x"26D2" => data <= "00000";
                when x"26D3" => data <= "10001";
                when x"26D4" => data <= "00110";
                when x"26D5" => data <= "00000";
                when x"26D6" => data <= "00000";
                when x"26D7" => data <= "00000";
                when x"26D8" => data <= "00000";
                when x"26D9" => data <= "00001";
                when x"26DA" => data <= "10111";
                when x"26DB" => data <= "00000";
                when x"26DC" => data <= "11010";
                when x"26DD" => data <= "00000";
                when x"26DE" => data <= "00110";
                when x"26DF" => data <= "10011";
                when x"26E0" => data <= "00110";
                when x"26E1" => data <= "00000";
                when x"26E2" => data <= "10011";
                when x"26E3" => data <= "00000";
                when x"26E4" => data <= "11011";
                when x"26E5" => data <= "00110";
                when x"26E6" => data <= "00110";
                when x"26E7" => data <= "00000";
                when x"26E8" => data <= "00000";
                when x"26E9" => data <= "00000";
                when x"26EA" => data <= "00000";
                when x"26EB" => data <= "00110";
                when x"26EC" => data <= "00110";
                when x"26ED" => data <= "00000";
                when x"26EE" => data <= "00000";
                when x"26EF" => data <= "00110";
                when x"26F0" => data <= "00000";
                when x"26F1" => data <= "01011";
                when x"26F2" => data <= "00000";
                when x"26F3" => data <= "00110";
                when x"26F4" => data <= "00000";
                when x"26F5" => data <= "00000";
                when x"26F6" => data <= "00110";
                when x"26F7" => data <= "00000";
                when x"26F8" => data <= "00110";
                when x"26F9" => data <= "10101";
                when x"26FA" => data <= "11010";
                when x"26FB" => data <= "00000";
                when x"26FC" => data <= "00000";
                when x"26FD" => data <= "00000";
                when x"26FE" => data <= "00011";
                when x"26FF" => data <= "00000";
                when x"2700" => data <= "11110";
                when x"2701" => data <= "00110";
                when x"2702" => data <= "00000";
                when x"2703" => data <= "00000";
                when x"2704" => data <= "00000";
                when x"2705" => data <= "00000";
                when x"2706" => data <= "00000";
                when x"2707" => data <= "00000";
                when x"2708" => data <= "00110";
                when x"2709" => data <= "00110";
                when x"270A" => data <= "01101";
                when x"270B" => data <= "11100";
                when x"270C" => data <= "00000";
                when x"270D" => data <= "10111";
                when x"270E" => data <= "00110";
                when x"270F" => data <= "00000";
                when x"2710" => data <= "00000";
                when x"2711" => data <= "01110";
                when x"2712" => data <= "00110";
                when x"2713" => data <= "00000";
                when x"2714" => data <= "00110";
                when x"2715" => data <= "11011";
                when x"2716" => data <= "10011";
                when x"2717" => data <= "00000";
                when x"2718" => data <= "00110";
                when x"2719" => data <= "00110";
                when x"271A" => data <= "00110";
                when x"271B" => data <= "00110";
                when x"271C" => data <= "00110";
                when x"271D" => data <= "00000";
                when x"271E" => data <= "00110";
                when x"271F" => data <= "01011";
                when x"2720" => data <= "10011";
                when x"2721" => data <= "00110";
                when x"2722" => data <= "00110";
                when x"2723" => data <= "00000";
                when x"2724" => data <= "00110";
                when x"2725" => data <= "00001";
                when x"2726" => data <= "00110";
                when x"2727" => data <= "00001";
                when x"2728" => data <= "11110";
                when x"2729" => data <= "00000";
                when x"272A" => data <= "00110";
                when x"272B" => data <= "00000";
                when x"272C" => data <= "00000";
                when x"272D" => data <= "00000";
                when x"272E" => data <= "01100";
                when x"272F" => data <= "00000";
                when x"2730" => data <= "00000";
                when x"2731" => data <= "01010";
                when x"2732" => data <= "01011";
                when x"2733" => data <= "00110";
                when x"2734" => data <= "00110";
                when x"2735" => data <= "00110";
                when x"2736" => data <= "00000";
                when x"2737" => data <= "00001";
                when x"2738" => data <= "00000";
                when x"2739" => data <= "00110";
                when x"273A" => data <= "00000";
                when x"273B" => data <= "10110";
                when x"273C" => data <= "00110";
                when x"273D" => data <= "00110";
                when x"273E" => data <= "00111";
                when x"273F" => data <= "00000";
                when x"2740" => data <= "00110";
                when x"2741" => data <= "00000";
                when x"2742" => data <= "00110";
                when x"2743" => data <= "00000";
                when x"2744" => data <= "00000";
                when x"2745" => data <= "00000";
                when x"2746" => data <= "10010";
                when x"2747" => data <= "00110";
                when x"2748" => data <= "00110";
                when x"2749" => data <= "00110";
                when x"274A" => data <= "00110";
                when x"274B" => data <= "00110";
                when x"274C" => data <= "00000";
                when x"274D" => data <= "00000";
                when x"274E" => data <= "00000";
                when x"274F" => data <= "00110";
                when x"2750" => data <= "01011";
                when x"2751" => data <= "00001";
                when x"2752" => data <= "00000";
                when x"2753" => data <= "00110";
                when x"2754" => data <= "01100";
                when x"2755" => data <= "00110";
                when x"2756" => data <= "00000";
                when x"2757" => data <= "00110";
                when x"2758" => data <= "00000";
                when x"2759" => data <= "00000";
                when x"275A" => data <= "00000";
                when x"275B" => data <= "00000";
                when x"275C" => data <= "00110";
                when x"275D" => data <= "00110";
                when x"275E" => data <= "00000";
                when x"275F" => data <= "00000";
                when x"2760" => data <= "00000";
                when x"2761" => data <= "00000";
                when x"2762" => data <= "00110";
                when x"2763" => data <= "00000";
                when x"2764" => data <= "00000";
                when x"2765" => data <= "00110";
                when x"2766" => data <= "00000";
                when x"2767" => data <= "01110";
                when x"2768" => data <= "10111";
                when x"2769" => data <= "10011";
                when x"276A" => data <= "00110";
                when x"276B" => data <= "11111";
                when x"276C" => data <= "11011";
                when x"276D" => data <= "00000";
                when x"276E" => data <= "00000";
                when x"276F" => data <= "00000";
                when x"2770" => data <= "00000";
                when x"2771" => data <= "00110";
                when x"2772" => data <= "00000";
                when x"2773" => data <= "00110";
                when x"2774" => data <= "00110";
                when x"2775" => data <= "00110";
                when x"2776" => data <= "00000";
                when x"2777" => data <= "00000";
                when x"2778" => data <= "00100";
                when x"2779" => data <= "00110";
                when x"277A" => data <= "00000";
                when x"277B" => data <= "00110";
                when x"277C" => data <= "00111";
                when x"277D" => data <= "00110";
                when x"277E" => data <= "00110";
                when x"277F" => data <= "00110";
                when x"2780" => data <= "00000";
                when x"2781" => data <= "00000";
                when x"2782" => data <= "00110";
                when x"2783" => data <= "00000";
                when x"2784" => data <= "01011";
                when x"2785" => data <= "00110";
                when x"2786" => data <= "00000";
                when x"2787" => data <= "00000";
                when x"2788" => data <= "00000";
                when x"2789" => data <= "00110";
                when x"278A" => data <= "00000";
                when x"278B" => data <= "10101";
                when x"278C" => data <= "00110";
                when x"278D" => data <= "00110";
                when x"278E" => data <= "00000";
                when x"278F" => data <= "00110";
                when x"2790" => data <= "00110";
                when x"2791" => data <= "10100";
                when x"2792" => data <= "11101";
                when x"2793" => data <= "00000";
                when x"2794" => data <= "00000";
                when x"2795" => data <= "00110";
                when x"2796" => data <= "00110";
                when x"2797" => data <= "00110";
                when x"2798" => data <= "00110";
                when x"2799" => data <= "11001";
                when x"279A" => data <= "00000";
                when x"279B" => data <= "00000";
                when x"279C" => data <= "10011";
                when x"279D" => data <= "00000";
                when x"279E" => data <= "00000";
                when x"279F" => data <= "01101";
                when x"27A0" => data <= "11001";
                when x"27A1" => data <= "00000";
                when x"27A2" => data <= "00110";
                when x"27A3" => data <= "00110";
                when x"27A4" => data <= "00110";
                when x"27A5" => data <= "00110";
                when x"27A6" => data <= "00110";
                when x"27A7" => data <= "00000";
                when x"27A8" => data <= "00101";
                when x"27A9" => data <= "00000";
                when x"27AA" => data <= "00110";
                when x"27AB" => data <= "00110";
                when x"27AC" => data <= "00110";
                when x"27AD" => data <= "00110";
                when x"27AE" => data <= "01001";
                when x"27AF" => data <= "00110";
                when x"27B0" => data <= "00110";
                when x"27B1" => data <= "00110";
                when x"27B2" => data <= "00110";
                when x"27B3" => data <= "00110";
                when x"27B4" => data <= "00000";
                when x"27B5" => data <= "00000";
                when x"27B6" => data <= "00110";
                when x"27B7" => data <= "00110";
                when x"27B8" => data <= "00110";
                when x"27B9" => data <= "00110";
                when x"27BA" => data <= "00110";
                when x"27BB" => data <= "00000";
                when x"27BC" => data <= "00010";
                when x"27BD" => data <= "00100";
                when x"27BE" => data <= "00110";
                when x"27BF" => data <= "00110";
                when x"27C0" => data <= "00110";
                when x"27C1" => data <= "00000";
                when x"27C2" => data <= "00110";
                when x"27C3" => data <= "01111";
                when x"27C4" => data <= "00010";
                when x"27C5" => data <= "00000";
                when x"27C6" => data <= "00000";
                when x"27C7" => data <= "00110";
                when x"27C8" => data <= "00110";
                when x"27C9" => data <= "00110";
                when x"27CA" => data <= "00000";
                when x"27CB" => data <= "00000";
                when x"27CC" => data <= "00000";
                when x"27CD" => data <= "01011";
                when x"27CE" => data <= "00110";
                when x"27CF" => data <= "00110";
                when x"27D0" => data <= "00110";
                when x"27D1" => data <= "00110";
                when x"27D2" => data <= "10011";
                when x"27D3" => data <= "00110";
                when x"27D4" => data <= "00110";
                when x"27D5" => data <= "00110";
                when x"27D6" => data <= "00000";
                when x"27D7" => data <= "00000";
                when x"27D8" => data <= "00000";
                when x"27D9" => data <= "00110";
                when x"27DA" => data <= "00110";
                when x"27DB" => data <= "00000";
                when x"27DC" => data <= "00000";
                when x"27DD" => data <= "00000";
                when x"27DE" => data <= "00000";
                when x"27DF" => data <= "00000";
                when x"27E0" => data <= "01011";
                when x"27E1" => data <= "00000";
                when x"27E2" => data <= "00000";
                when x"27E3" => data <= "00110";
                when x"27E4" => data <= "00110";
                when x"27E5" => data <= "00110";
                when x"27E6" => data <= "00101";
                when x"27E7" => data <= "00110";
                when x"27E8" => data <= "00000";
                when x"27E9" => data <= "00110";
                when x"27EA" => data <= "00001";
                when x"27EB" => data <= "00000";
                when x"27EC" => data <= "11101";
                when x"27ED" => data <= "00110";
                when x"27EE" => data <= "01011";
                when x"27EF" => data <= "10100";
                when x"27F0" => data <= "01001";
                when x"27F1" => data <= "00000";
                when x"27F2" => data <= "00110";
                when x"27F3" => data <= "01010";
                when x"27F4" => data <= "00000";
                when x"27F5" => data <= "00000";
                when x"27F6" => data <= "00000";
                when x"27F7" => data <= "10011";
                when x"27F8" => data <= "11011";
                when x"27F9" => data <= "00110";
                when x"27FA" => data <= "01100";
                when x"27FB" => data <= "00000";
                when x"27FC" => data <= "00110";
                when x"27FD" => data <= "00110";
                when x"27FE" => data <= "00110";
                when x"27FF" => data <= "10101";
                when others => data <= (others => '0');
            end case;
        end if;
    end process;
end Behavioral;




----------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


entity reading_normal is
    generic (
        dimension_size     : integer := 1024;   -- dimension size 
        dimension_WIDTH    : integer := 10;     -- log2 dimension size 
        class_size    : integer := 10;     -- number of classes
        ECC_WIDTH          : integer := 8       -- bit-width of ECC_code 
    );
	port (
	clk                     : in std_logic;
    rst                     : in std_logic;
	din 					: in std_logic_vector(dimension_size-1 downto 0);
    count_reg               : in std_logic_vector(dimension_WIDTH-1 downto 0);
    dout                    : out std_logic_vector(dimension_WIDTH-1 downto 0)
	);	
end entity;

architecture behavior of reading_normal is

    -- Array types
    type CHV_memory_array is array (0 to dimension_size-1) of std_logic_vector(class_size-1 downto 0);
    type countingCheck is array (0 to dimension_WIDTH-1) of std_logic_vector(dimension_WIDTH-1 downto 0);

    -- Signals
    signal CHV_memory               : CHV_memory_array;
    signal CHV_memory_out : std_logic_vector(class_size-1 downto 0);
    signal corrected_CHV_memory_out : std_logic_vector(class_size-1 downto 0);

    signal count_sim               : countingCheck;
    signal double_error    : std_logic;

    -- File I/O
    
    signal en_pops_regular         : std_logic_vector(class_size-1 downto 0);
    
    signal LFSRasHVCheck           : std_logic;
    signal LFSR_suffleAsHVCheck    : std_logic;

	signal ECC_out             : std_logic_vector(5-1 downto 0);
    
begin

    CHVMem: entity work.CHV_mem_10000
    port map(
    clk  => clk,
    address => count_reg,
    data => CHV_memory_out
    );
    
	ECCuut: entity work.ECC_vhdl_module
    generic map(
        C  => class_size,
        ECC_bit => 5   )
    port map(
        d => CHV_memory_out,
        p => ECC_out,
        double_error => double_error,
        dcw   => corrected_CHV_memory_out
    );
    
	ECCuutMem: entity work.ECC_CHV_img_10000
    port map(
    clk  => clk,
    address => count_reg,
    data => ECC_out
    );

    LFSRasHVCheck  <= din(to_integer(unsigned(count_reg)));

    en_regular_pops: for k in 0 to class_size-1 generate
        en_pops_regular(k) <= corrected_CHV_memory_out(k) xor LFSRasHVCheck;
    end generate;

    -- Counters for regular
    class_counter: for k in 0 to class_size-1 generate
        simcounter: entity work.popCount 
            generic map(lenPop => dimension_WIDTH)
            port map(
                clk  => clk,
                rst  => rst,
                en   => en_pops_regular(k),
                dout => count_sim(k)
            );
    end generate;
	
	dout <= std_logic_vector(unsigned(count_sim(0)) + unsigned(count_sim(1)) + unsigned(count_sim(2)) + unsigned(count_sim(3)) + unsigned(count_sim(4)) + unsigned(count_sim(5)) + unsigned(count_sim(6)) + unsigned(count_sim(7)) + unsigned(count_sim(8)) + unsigned(count_sim(9)));
end architecture;



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity top_module_for_normal_ECC_10000 is
    generic (
        dimension_size     : integer := 10240;   -- dimension size 
        dimension_WIDTH    : integer := 14;     -- log2 dimension size 
        dimension_segmentation    : integer := 1280;     -- genrate input
        class_size    : integer := 10;     -- number of classes
        ECC_WIDTH          : integer := 5       -- bit-width of ECC_code 
    );
    port (
	clk                     : in std_logic;
    rst                     : in std_logic;
    pop_en                  : in std_logic;
	din 					: in std_logic_vector((dimension_size/dimension_segmentation)-1 downto 0);
      count_sim     :out std_logic_vector(dimension_WIDTH-1 downto 0)
	);	
end entity;

architecture behavior of top_module_for_normal_ECC_10000 is

signal realdin 					:  std_logic_vector((dimension_size)-1 downto 0);

type index_array is array (0 to dimension_size-1) of std_logic_vector(dimension_WIDTH-1 downto 0);
    
signal index_memory               : index_array;
signal count_reg               :  std_logic_vector(dimension_WIDTH-1 downto 0);
       
begin

    input_gen: for k in 0 to dimension_segmentation-1 generate
        realdin((dimension_size/dimension_segmentation)*(k+1)-1 downto (dimension_size/dimension_segmentation)*k) <= din;
    end generate;
    
    
    ECCuutMem: entity work.reading_normal 
	generic map(
		dimension_size  => dimension_size,
        dimension_WIDTH  => dimension_WIDTH,
        class_size  =>  class_size,
        ECC_WIDTH => ECC_WIDTH)
	port map(
		clk  => clk,
		rst  => rst,
		din  => realdin,
	    count_reg 		=> count_reg,
		dout  => count_sim
		);

    -- Count_reg counter
    counter: entity work.popCount 
        generic map(lenPop => dimension_WIDTH)
        port map(
            clk  => clk,
            rst  => rst,
            en   => pop_en,
            dout => count_reg
        );

end architecture;
